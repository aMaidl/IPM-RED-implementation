/****************************************************************************

 * roundAES.v

 ****************************************************************************/



/**

 * Module: roundAES

 * 

 * TODO: Add module documentation

 */
module roundAES #(parameter v = 3) (
	input  clk,
	input  rst,
	input  en,
	input [16*(v*8)-1:0] plaintext,
	input [16*(v*8)-1:0] round_ks,
	input [(v*8)-1:0] L,
	input [(v*v*8)-1:0] L_hat,
	input [2*80-1:0] RNG_seed,
	output reg can_supply_last,
	output [3:0] current_round,
	output [16*(v*8)-1:0] ciphertext,
	output reg is_busy
);


    parameter BRAM_mul = 3'b000;
    parameter BRAM_add = 3'b001;
    parameter BRAM_sq = 3'b010;
    parameter BRAM_mc = 3'b011;
    parameter BRAM_PT = 3'b100;
    parameter BRAM_KS = 3'b101;
    parameter BRAM_mask = 3'b110;
    parameter BRAM_DEFAULT = 3'b111;


	wire [(v*v*8)-2:0] IPMMult_rand;
	wire [(v-1)*8-1:0] IPMMask_rand;
	wire RNGisReady;

	reg RNGenable;
	reg RNGreseed;
	reg RNGisInit = 0;

    RNG_Trivium64 #(.instances(2)) RNG_Trivium64 (
        .clk(clk),
        .enable(en),
        .reseed(RNGreseed),
        .seed(RNG_seed),
        .isReady(RNGisReady),
        .random({IPMMult_rand, IPMMask_rand})
    );


    reg [16*(v*8)-1:0] round_pt;

	//==============================
	// wires :
	//==============================


	wire  [v*8-1:0] IPMSquare_Z;
	wire [v*8-1:0] IPMSquare_P;
	wire  [v*8-1:0] IPMMult_Z;
	wire  [v*8-1:0] IPMMult_Z_;
	wire [v*8-1:0] IPMMult_P;
	wire  [v*8-1:0] IPMAdd_Z;
	wire  [v*8-1:0] IPMAdd_Z_;
	wire [v*8-1:0] IPMAdd_P;
	wire [v*8-1:0] IPMMask_R;
	wire  [v*8-1:0] IPMMultConst_Z;
	reg  [8-1:0] IPMMultConst_const;
	wire [v*8-1:0] IPMMultConst_P;


	reg  [10-1:0] state;
	reg  [3:0] round_count;
	assign current_round = round_count;

	//==============================
	// IO :
	//==============================
	assign ciphertext = round_pt;

	//==============================
	// modules :
	//==============================
	IPSquare #(.v(v)) IPSquare(
		.R(IPMSquare_Z),
		.L(L),
		.T(IPMSquare_P)
	);

	IPMult #(.v(v)) IPMult(
		.rand(IPMMult_rand),
		.R(IPMMult_Z),
		.Q(IPMMult_Z_),
		.L_hat(L_hat),
		.T(IPMMult_P)
	);

	IPAdd #(.v(v)) IPAdd(
		.R(IPMAdd_Z),
		.Q(IPMAdd_Z_),
		.T(IPMAdd_P)
	);

	IPMask #(.v(v)) IPMask(
		.rand(IPMMask_rand),
		.S(8'h63),
		.L(L),
		.R(IPMMask_R)
	);

	IPMultConst #(.v(v)) IPMultConst(
		.R(IPMMultConst_Z),
		.const(IPMMultConst_const),
		.T(IPMMultConst_P)
	);



	reg IPMAdd_BRAM_en;
	reg IPMMult_BRAM_en;
	reg IPMMultConst_BRAM_en;
	reg IPMSquare_BRAM_en;
	reg [4:0] IPMAdd_addr_w;
	reg [4:0] IPMMult_addr_w;
	reg [4:0] IPMMultConst_addr_w;
	reg [4:0] IPMSquare_addr_w;

    reg [4:0] IPMAdd_Z_addr_r;
    reg [4:0] IPMAdd_Z__addr_r;
    reg [4:0] IPMMult_Z_addr_r;
    reg [4:0] IPMMult_Z__addr_r;
    reg [4:0] IPMMultConst_Z_addr_r;
    reg [4:0] IPMSquare_Z_addr_r;

    reg [2:0] IPMAdd_Z_addr_r_BRAM;
    reg [2:0] IPMAdd_Z__addr_r_BRAM;
    reg [2:0] IPMMult_Z_addr_r_BRAM;
    reg [2:0] IPMMult_Z__addr_r_BRAM;
    reg [2:0] IPMMultConst_Z_addr_r_BRAM;
    reg [2:0] IPMSquare_Z_addr_r_BRAM;

    Bank #(.addr_bits(5), .debug(1)) Bank (
         .DEBUG_STATE(state),
         .clk(clk),
         .en(en),
         .plaintext(round_pt),
         .round_ks(round_ks),
         .add_en(IPMAdd_BRAM_en),
         .mul_en(IPMMult_BRAM_en),
         .mc_en(IPMMultConst_BRAM_en),
         .sq_en(IPMSquare_BRAM_en),
         .add_addr_w(IPMAdd_addr_w),
         .mul_addr_w(IPMMult_addr_w),
         .mc_addr_w(IPMMultConst_addr_w),
         .sq_addr_w(IPMSquare_addr_w),
         .add_val_w(IPMAdd_P),
         .mul_val_w(IPMMult_P),
         .mc_val_w(IPMMultConst_P),
         .sq_val_w(IPMSquare_P),
         .mask_val_w(IPMMask_R),
         .add0_addr_r(IPMAdd_Z_addr_r),
         .add1_addr_r(IPMAdd_Z__addr_r),
         .mul0_addr_r(IPMMult_Z_addr_r),
         .mul1_addr_r(IPMMult_Z__addr_r),
         .mc_addr_r(IPMMultConst_Z_addr_r),
         .sq_addr_r(IPMSquare_Z_addr_r),
         .add0_r_BRAM(IPMAdd_Z_addr_r_BRAM),
         .add1_r_BRAM(IPMAdd_Z__addr_r_BRAM),
         .mul0_r_BRAM(IPMMult_Z_addr_r_BRAM),
         .mul1_r_BRAM(IPMMult_Z__addr_r_BRAM),
         .mc_r_BRAM(IPMMultConst_Z_addr_r_BRAM),
         .sq_r_BRAM(IPMSquare_Z_addr_r_BRAM),
         .add0_out(IPMAdd_Z),
         .add1_out(IPMAdd_Z_),
         .mul0_out(IPMMult_Z),
         .mul1_out(IPMMult_Z_),
         .mc_out(IPMMultConst_Z),
         .sq_out(IPMSquare_Z)
    );




	//==============================
	// control :
	//==============================


	wire is_last = (round_count == 10);
	always @(posedge clk) begin
		if (!rst) begin
			state <= 10'b1111111111;
			is_busy <= 1;
		end
		else begin
            if(!en) begin
                state <= 10'b1111111111;
					 is_busy <= 1;
            end else begin
                $display("=====================");
                $display("state       = %b (%d)", state, state);
                $display("round_count = %d", round_count);
                $display("L          = %h" , L);
                $display("L_hat      = %h" , L_hat);
                $display("rpt        = %h", round_pt);
                $display("round_ks   = %h", round_ks);
                //$display("r1          = %h", IPMMult_rand);
                //$display("r2          = %h", IPMAdd_rand);
                //$display("r3          = %h", IPMMask_rand);
                /*
                $display("(%d) +  um = %h", state, add_um);
                $display("(%d) *  um = %h", state, mul_um);
                $display("(%d) mc um = %h", state, mc_um);
                $display("(%d) sq um = %h", state, sq_um);
                */



                // these are important!!!
                IPMAdd_BRAM_en <= 0;
                IPMMult_BRAM_en <= 0;
                IPMMultConst_BRAM_en <= 0;
                IPMSquare_BRAM_en <= 0;
                IPMAdd_Z_addr_r_BRAM <= BRAM_DEFAULT;
                IPMAdd_Z__addr_r_BRAM <= BRAM_DEFAULT;
                IPMMult_Z_addr_r_BRAM <= BRAM_DEFAULT;
                IPMMult_Z__addr_r_BRAM <= BRAM_DEFAULT;
                IPMSquare_Z_addr_r_BRAM <= BRAM_DEFAULT;
                IPMMultConst_Z_addr_r_BRAM <= BRAM_DEFAULT;
                IPMMultConst_const <= 8'h0;
                // 0 address is not in use
                IPMSquare_addr_w <= 8'h0;
                IPMMult_addr_w <= 8'h0;
                IPMAdd_addr_w <= 8'h0;
                IPMMultConst_addr_w <= 8'h0;

                // FSM
                case(state)                    // reset RNG
                    10'b1111111111 : begin
                        can_supply_last <= 0;
                        RNGreseed <= 1;
                        RNGenable <= 1;
                        state <= 10'b1111111110;
                        round_count <= 1;
                        round_pt <= plaintext[1*16*v*8-1:0*16*v*8];
								is_busy <= 1;
                    end
                    // wait until RNG is ready
                    10'b1111111110 : begin
                        RNGreseed <= 0;
                        if (RNGisReady) begin
                            state <= 10'b0000000000;
                        end else begin
                            state <= 10'b1111111110;
                        end
                    end
                    // rounds 1-9 start here
                   10'b0000000000 : begin
                   	state <= 10'b0000000001;
                   	IPMAdd_Z_addr_r <= 5'h10; // addr of byte F
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h10; // addr of byte F
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   end
                   10'b0000000001 : begin
                   	state <= 10'b0000000010;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hF; // addr of byte E
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hF; // addr of byte E
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMSquare_Z_addr_r <= 5'h11;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000000010 : begin
						 
                   	state <= 10'b0000000011;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hE; // addr of byte D
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hE; // addr of byte D
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h11;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000000011 : begin
						 
                   	
                   	state <= 10'b0000000100;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hD; // addr of byte C
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hD; // addr of byte C
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMult_addr_w <= 5'h15;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hA;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h15;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000000100 : begin
						 
                   	
                   	state <= 10'b0000000101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hC; // addr of byte B
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hC; // addr of byte B
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMult_addr_w <= 5'h19;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h11;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000000101 : begin
						 
                   	
                   	state <= 10'b0000000110;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hB; // addr of byte A
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hB; // addr of byte A
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMMult_addr_w <= 5'h16;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hE;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000000110 : begin
						 
                   	
                   	
                   	state <= 10'b0000000111;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hA; // addr of byte 9
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hA; // addr of byte 9
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMult_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h15;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h19;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000000111 : begin
						 
                   	
                   	
                   	state <= 10'b0000001000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h9; // addr of byte 8
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h9; // addr of byte 8
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h16;
                   	IPMMult_addr_w <= 5'h15;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hA;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000001000 : begin
						 
                   	
                   	
                   	state <= 10'b0000001001;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h8; // addr of byte 7
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h8; // addr of byte 7
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMult_addr_w <= 5'h13;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h3;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h11;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000001001 : begin
						 
                   	
                   	
                   	state <= 10'b0000001010;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h7; // addr of byte 6
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h7; // addr of byte 6
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMult_addr_w <= 5'h9;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h11;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000001010 : begin
						 
                   	
                   	
                   	state <= 10'b0000001011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h6; // addr of byte 5
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h6; // addr of byte 5
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h13;
                   	IPMMult_addr_w <= 5'h1C;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hE;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000001011 : begin
						 
                   	
                   	
                   	state <= 10'b0000001100;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h5; // addr of byte 4
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h5; // addr of byte 4
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMult_addr_w <= 5'hE;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMMult_Z_addr_r <= 5'h3;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h15;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000001100 : begin
						 
                   	
                   	
                   	state <= 10'b0000001101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h4; // addr of byte 3
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h4; // addr of byte 3
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMult_addr_w <= 5'h15;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000001101 : begin
						 
                   	
                   	
                   	state <= 10'b0000001110;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h3; // addr of byte 2
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h3; // addr of byte 2
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h19;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h16;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000001110 : begin
						 
                   	
                   	
                   	state <= 10'b0000001111;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h2; // addr of byte 1
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h2; // addr of byte 1
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMult_addr_w <= 5'h19;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h16;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000001111 : begin
						 
                   	
                   	
                   	state <= 10'b0000010000;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h1; // addr of byte 0
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h1; // addr of byte 0
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h1B;
                   	IPMMult_addr_w <= 5'h12;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hA;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000010000 : begin
						 
                   	
                   	
                   	state <= 10'b0000010001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h14;
                   	IPMMult_addr_w <= 5'h18;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h3;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000010001 : begin
						 
                   	
                   	
                   	state <= 10'b0000010010;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hF;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000010010 : begin
                   	state <= 10'b0000010011;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h17;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h8;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h1C;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000010011 : begin
                   	state <= 10'b0000010100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h11;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h13;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000010100 : begin
                   	state <= 10'b0000010101;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hC;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h13;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000010101 : begin
                   	state <= 10'b0000010110;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h1B;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hE;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000010110 : begin
                   	state <= 10'b0000010111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h1A;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMSquare_Z_addr_r <= 5'h15;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000010111 : begin
                   	state <= 10'b0000011000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000011000 : begin
                   	state <= 10'b0000011001;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMMult_Z_addr_r <= 5'hA;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h2;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000011001 : begin
                   	state <= 10'b0000011010;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h14;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMMult_Z_addr_r <= 5'hA;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h8;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h19;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000011010 : begin
                   	state <= 10'b0000011011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h19;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000011011 : begin
                   	state <= 10'b0000011100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h7;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h12;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000011100 : begin
                   	state <= 10'b0000011101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h11;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h16;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h1B;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000011101 : begin
                   	state <= 10'b0000011110;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1B;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000011110 : begin
                   	state <= 10'b0000011111;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hD;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h9;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h18;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000011111 : begin
                   	state <= 10'b0000100000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h9;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hA;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h14;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000100000 : begin
                   	state <= 10'b0000100001;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h2;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h14;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h17;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000100001 : begin
                   	state <= 10'b0000100010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hF;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hF;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000100010 : begin
                   	state <= 10'b0000100011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000100011 : begin
                   	state <= 10'b0000100100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1C;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h1B;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000100100 : begin
                   	state <= 10'b0000100101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h1C;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h13;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000100101 : begin
                   	state <= 10'b0000100110;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMMult_Z_addr_r <= 5'h3;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h16;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h1A;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000100110 : begin
                   	state <= 10'b0000100111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h16;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMMult_Z_addr_r <= 5'h3;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hE;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h16;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000100111 : begin
                   	state <= 10'b0000101000;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMult_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h15;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h14;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000101000 : begin
                   	state <= 10'b0000101001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMult_addr_w <= 5'h15;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h2;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000101001 : begin
                   	state <= 10'b0000101010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h5;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMSquare_Z_addr_r <= 5'h19;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000101010 : begin
                   	state <= 10'b0000101011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMMult_Z_addr_r <= 5'hD;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h8;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000101011 : begin
                   	state <= 10'b0000101100;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h12;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h11;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000101100 : begin
                   	state <= 10'b0000101101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h12;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h7;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000101101 : begin
                   	state <= 10'b0000101110;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMMult_Z_addr_r <= 5'h4;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1B;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000101110 : begin
                   	state <= 10'b0000101111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h9;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000101111 : begin
                   	state <= 10'b0000110000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h18;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000110000 : begin
                   	state <= 10'b0000110001;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h18;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h17;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000110001 : begin
                   	state <= 10'b0000110010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h17;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h14;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000110010 : begin
                   	state <= 10'b0000110011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMSquare_Z_addr_r <= 5'h1C;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000110011 : begin
                   	state <= 10'b0000110100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000110100 : begin
                   	state <= 10'b0000110101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1B;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h16;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000110101 : begin
                   	state <= 10'b0000110110;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h16;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000110110 : begin
                   	state <= 10'b0000110111;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'h3;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1A;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h15;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000110111 : begin
                   	state <= 10'b0000111000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMult_addr_w <= 5'h15;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111000 : begin
                   	state <= 10'b0000111001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h14;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111001 : begin
                   	state <= 10'b0000111010;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h14;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMMult_Z_addr_r <= 5'hA;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h13;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111010 : begin
                   	state <= 10'b0000111011;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h13;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMMult_Z_addr_r <= 5'hD;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h19;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h13;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h12;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000111011 : begin
                   	state <= 10'b0000111100;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMult_addr_w <= 5'h12;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111100 : begin
                   	state <= 10'b0000111101;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h14;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h11;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111101 : begin
                   	state <= 10'b0000111110;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h11;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMMult_Z_addr_r <= 5'h4;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hD;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111110 : begin
                   	state <= 10'b0000111111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hD;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMSquare_Z_addr_r <= 5'h18;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000111111 : begin
                   	state <= 10'b0001000000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMSquare_Z_addr_r <= 5'h17;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001000000 : begin
                   	state <= 10'b0001000001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001000001 : begin
                   	state <= 10'b0001000010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hF;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001000010 : begin
                   	state <= 10'b0001000011;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hF;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMMult_Z_addr_r <= 5'hB;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hE;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001000011 : begin
                   	state <= 10'b0001000100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hE;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001000100 : begin
                   	state <= 10'b0001000101;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h16;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001000101 : begin
                   	state <= 10'b0001000110;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1B;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001000110 : begin
                   	state <= 10'b0001000111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMSquare_Z_addr_r <= 5'h15;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001000111 : begin
                   	state <= 10'b0001001000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMSquare_Z_addr_r <= 5'h14;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001001000 : begin
                   	state <= 10'b0001001001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMSquare_Z_addr_r <= 5'h13;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001001001 : begin
                   	state <= 10'b0001001010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001001010 : begin
                   	state <= 10'b0001001011;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h14;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h12;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001001011 : begin
                   	state <= 10'b0001001100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h14;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMSquare_Z_addr_r <= 5'h11;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001001100 : begin
                   	state <= 10'b0001001101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001001101 : begin
                   	state <= 10'b0001001110;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMMult_Z_addr_r <= 5'h9;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h10;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001001110 : begin
                   	state <= 10'b0001001111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hD;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001001111 : begin
                   	state <= 10'b0001010000;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010000 : begin
                   	state <= 10'b0001010001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001010001 : begin
                   	state <= 10'b0001010010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001010010 : begin
                   	state <= 10'b0001010011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010011 : begin
                   	state <= 10'b0001010100;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1B;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hC;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010100 : begin
                   	state <= 10'b0001010101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1B;
                   	IPMMult_addr_w <= 5'hC;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010101 : begin
                   	state <= 10'b0001010110;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010110 : begin
                   	state <= 10'b0001010111;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMult_Z_addr_r <= 5'h3;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h7;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010111 : begin
                   	state <= 10'b0001011000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMult_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011000 : begin
                   	state <= 10'b0001011001;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011001 : begin
                   	state <= 10'b0001011010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011010 : begin
                   	state <= 10'b0001011011;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h14;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'hD;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hA;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011011 : begin
                   	state <= 10'b0001011100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h14;
                   	IPMMult_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011100 : begin
                   	state <= 10'b0001011101;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001011101 : begin
                   	state <= 10'b0001011110;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h13;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011110 : begin
                   	state <= 10'b0001011111;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011111 : begin
                   	state <= 10'b0001100000;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMMult_Z_addr_r <= 5'h4;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h2;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100000 : begin
                   	state <= 10'b0001100001;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h2;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h8;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100001 : begin
                   	state <= 10'b0001100010;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMult_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100010 : begin
                   	state <= 10'b0001100011;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100011 : begin
                   	state <= 10'b0001100100;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1B;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001100100 : begin
                   	state <= 10'b0001100101;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1B;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100101 : begin
                   	state <= 10'b0001100110;
                   	IPMMultConst_const <= 8'h5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'hB;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hB;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001100110 : begin
                   	state <= 10'b0001100111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMult_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100111 : begin
                   	state <= 10'b0001101000;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h6;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101000 : begin
                   	state <= 10'b0001101001;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMult_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMult_Z_addr_r <= 5'hA;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h5;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101001 : begin
                   	state <= 10'b0001101010;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'h16;
                   	IPMMult_addr_w <= 5'h5;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001101010 : begin
                   	state <= 10'b0001101011;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h14;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101011 : begin
                   	state <= 10'b0001101100;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'h14;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMult_Z_addr_r <= 5'h6;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h4;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101100 : begin
                   	state <= 10'b0001101101;
                   	IPMMultConst_const <= 8'h5;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMMult_addr_w <= 5'h4;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h13;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'h8;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h3;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101101 : begin
                   	state <= 10'b0001101110;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'h13;
                   	IPMMult_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101110 : begin
                   	state <= 10'b0001101111;
                   	IPMMultConst_const <= 8'h9;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'h9;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h9;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001101111 : begin
                   	state <= 10'b0001110000;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMult_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001110000 : begin
                   	state <= 10'b0001110001;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1C;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001110001 : begin
                   	state <= 10'b0001110010;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMult_Z_addr_r <= 5'h7;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001110010 : begin
                   	state <= 10'b0001110011;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h15;
                   	IPMMult_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001110011 : begin
                   	state <= 10'b0001110100;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1B;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001110100 : begin
                   	state <= 10'b0001110101;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'h1B;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001110101 : begin
                   	state <= 10'b0001110110;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001110110 : begin
                   	state <= 10'b0001110111;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001110111 : begin
                   	state <= 10'b0001111000;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001111000 : begin
                   	state <= 10'b0001111001;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h16;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001111001 : begin
                   	state <= 10'b0001111010;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h16;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001111010 : begin
                   	state <= 10'b0001111011;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h14;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001111011 : begin
                   	state <= 10'b0001111100;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h14;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001111100 : begin
                   	state <= 10'b0001111101;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h13;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001111101 : begin
                   	state <= 10'b0001111110;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h13;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001111110 : begin
                   	state <= 10'b0001111111;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001111111 : begin
                   	state <= 10'b0010000000;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1C;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000000 : begin
                   	state <= 10'b0010000001;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1C;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000001 : begin
                   	state <= 10'b0010000010;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h15;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0010000010 : begin
                   	state <= 10'b0010000011;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h15;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000011 : begin
                   	state <= 10'b0010000100;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000100 : begin
                   	state <= 10'b0010000101;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1B;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000101 : begin
                   	state <= 10'b0010000110;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1B;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000110 : begin
                   	state <= 10'b0010000111;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000111 : begin
                   	state <= 10'b0010001000;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001000 : begin
                   	state <= 10'b0010001001;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h16;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001001 : begin
                   	state <= 10'b0010001010;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h16;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001010 : begin
                   	state <= 10'b0010001011;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h14;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001011 : begin
                   	state <= 10'b0010001100;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h14;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001100 : begin
                   	state <= 10'b0010001101;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h13;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001101 : begin
                   	state <= 10'b0010001110;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h13;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001110 : begin
                   	state <= 10'b0010001111;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001111 : begin
                   	state <= 10'b0010010000;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1C;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010000 : begin
                   	state <= 10'b0010010001;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1C;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010001 : begin
                   	state <= 10'b0010010010;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h15;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010010 : begin
                   	state <= 10'b0010010011;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h15;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010011 : begin
                   	state <= 10'b0010010100;
                   	IPMMultConst_const <= 8'h9;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1B;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010100 : begin
                   	state <= 10'b0010010101;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1B;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010101 : begin
                   	state <= 10'b0010010110;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010110 : begin
                   	state <= 10'b0010010111;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010111 : begin
                   	state <= 10'b0010011000;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011000 : begin
                   	state <= 10'b0010011001;
                   	IPMMultConst_const <= 8'h2;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h16;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011001 : begin
                   	state <= 10'b0010011010;
                   	IPMMultConst_const <= 8'h3;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h16;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'hF;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h14;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011010 : begin
                   	state <= 10'b0010011011;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h14;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011011 : begin
                   	state <= 10'b0010011100;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011100 : begin
                   	state <= 10'b0010011101;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h13;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011101 : begin
                   	state <= 10'b0010011110;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h13;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011110 : begin
                   	state <= 10'b0010011111;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011111 : begin
                   	state <= 10'b0010100000;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1C;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100000 : begin
                   	state <= 10'b0010100001;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1C;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100001 : begin
                   	state <= 10'b0010100010;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'hE;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h1B;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100010 : begin
                   	state <= 10'b0010100011;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1B;
                   	IPMMultConst_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h15;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100011 : begin
                   	state <= 10'b0010100100;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h15;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'hB;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100100 : begin
                   	state <= 10'b0010100101;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100101 : begin
                   	state <= 10'b0010100110;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'hB;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100110 : begin
                   	state <= 10'b0010100111;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100111 : begin
                   	state <= 10'b0010101000;
                   	IPMMultConst_const <= 8'h25;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z__addr_r <= 5'hB;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h16;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101000 : begin
                   	state <= 10'b0010101001;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h16;
                   	IPMMultConst_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101001 : begin
                   	state <= 10'b0010101010;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'hB;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h14;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101010 : begin
                   	state <= 10'b0010101011;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h14;
                   	IPMMultConst_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101011 : begin
                   	state <= 10'b0010101100;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'hB;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h13;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h14;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101100 : begin
                   	state <= 10'b0010101101;
                   	IPMMultConst_const <= 8'h2;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h13;
                   	IPMMultConst_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'hD;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h14;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101101 : begin
                   	state <= 10'b0010101110;
                   	IPMMultConst_const <= 8'h3;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101110 : begin
                   	state <= 10'b0010101111;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1C;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101111 : begin
                   	state <= 10'b0010110000;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1C;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110000 : begin
                   	state <= 10'b0010110001;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h15;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110001 : begin
                   	state <= 10'b0010110010;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h15;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110010 : begin
                   	state <= 10'b0010110011;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1B;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110011 : begin
                   	state <= 10'b0010110100;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1B;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'hC;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1B;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110100 : begin
                   	state <= 10'b0010110101;
                   	IPMMultConst_const <= 8'h2;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'hE;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'hB;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1B;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110101 : begin
                   	state <= 10'b0010110110;
                   	IPMMultConst_const <= 8'h3;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h2;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110110 : begin
                   	state <= 10'b0010110111;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h16;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110111 : begin
                   	state <= 10'b0010111000;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h16;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h13;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111000 : begin
                   	state <= 10'b0010111001;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h13;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111001 : begin
                   	state <= 10'b0010111010;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111010 : begin
                   	state <= 10'b0010111011;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111011 : begin
                   	state <= 10'b0010111100;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111100 : begin
                   	state <= 10'b0010111101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h9;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111101 : begin
                   	state <= 10'b0010111110;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1C;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111110 : begin
                   	state <= 10'b0010111111;
                   	IPMMultConst_const <= 8'h2;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1C;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h8;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111111 : begin
                   	state <= 10'b0011000000;
                   	IPMMultConst_const <= 8'h3;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'hF;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h15;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000000 : begin
                   	state <= 10'b0011000001;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h15;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000001 : begin
                   	state <= 10'b0011000010;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000010 : begin
                   	state <= 10'b0011000011;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h16;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000011 : begin
                   	state <= 10'b0011000100;
                   	IPMMultConst_const <= 8'h2;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h16;
                   	IPMMultConst_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000100 : begin
                   	state <= 10'b0011000101;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000101 : begin
                   	state <= 10'b0011000110;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h9;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h5;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000110 : begin
                   	state <= 10'b0011000111;
                   	IPMMultConst_const <= 8'h2;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMMultConst_addr_w <= 5'h11;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'hE;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000111 : begin
                   	state <= 10'b0011001000;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h4;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001000 : begin
                   	state <= 10'b0011001001;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h9;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h13;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001001 : begin
                   	state <= 10'b0011001010;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h13;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001010 : begin
                   	state <= 10'b0011001011;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h9;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h1C;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h13;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001011 : begin
                   	state <= 10'b0011001100;
                   	IPMMultConst_const <= 8'h2;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1C;
                   	IPMMultConst_addr_w <= 5'hD;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h13;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001100 : begin
                   	state <= 10'b0011001101;
                   	IPMMultConst_const <= 8'h3;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hC;
                   	IPMMultConst_addr_w <= 5'h11;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z__addr_r <= 5'hE;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001101 : begin
                   	state <= 10'b0011001110;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001110 : begin
                   	state <= 10'b0011001111;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h2;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h15;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001111 : begin
                   	state <= 10'b0011010000;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h15;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h9;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011010000 : begin
                   	state <= 10'b0011010001;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'h9;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011010001 : begin
                   	state <= 10'b0011010010;
                   	IPMMultConst_const <= 8'h2;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'h5;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h16;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011010010 : begin
                   	state <= 10'b0011010011;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h16;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011010011 : begin
                   	state <= 10'b0011010100;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'hE;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011010100 : begin
                   	state <= 10'b0011010101;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h9;
                   	IPMMultConst_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'h1B;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011010101 : begin
                   	state <= 10'b0011010110;
                   	IPMMultConst_const <= 8'h2;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'h12;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011010110 : begin
                   	state <= 10'b0011010111;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMMultConst_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'h9;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011010111 : begin
                   	state <= 10'b0011011000;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h2;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h16;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011000 : begin
                   	state <= 10'b0011011001;
                   	IPMMultConst_const <= 8'h2;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1D;
                   	IPMMultConst_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h8;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h16;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h16;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011001 : begin
                   	state <= 10'b0011011010;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h8;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h16;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011010 : begin
                   	state <= 10'b0011011011;
                   	IPMMultConst_const <= 8'h2;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h16;
                   	IPMMultConst_addr_w <= 5'h8;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z__addr_r <= 5'h1B;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011011 : begin
                   	state <= 10'b0011011100;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1B;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1C;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h11;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011100 : begin
                   	state <= 10'b0011011101;
                   	IPMMultConst_const <= 8'h2;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1C;
                   	IPMMultConst_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'hE;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h15;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h11;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011101 : begin
                   	state <= 10'b0011011110;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h15;
                   	IPMMultConst_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'hD;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011110 : begin
                   	state <= 10'b0011011111;
                   	IPMMultConst_const <= 8'h2;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMMultConst_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h13;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011111 : begin
                   	state <= 10'b0011100000;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h11;
                   	IPMMultConst_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'h9;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1C;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100000 : begin
                   	state <= 10'b0011100001;
                   	IPMMultConst_const <= 8'h2;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h14;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1C;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100001 : begin
                   	state <= 10'b0011100010;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1A;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h15;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100010 : begin
                   	state <= 10'b0011100011;
                   	IPMMultConst_const <= 8'h2;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h15;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100011 : begin
                   	state <= 10'b0011100100;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h18;
                   	IPMMultConst_addr_w <= 5'h5;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z__addr_r <= 5'h8;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100100 : begin
                   	state <= 10'b0011100101;
                   	IPMMultConst_const <= 8'h2;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h1C;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100101 : begin
                   	state <= 10'b0011100110;
                   	IPMMultConst_const <= 8'h3;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1E;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h12;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1C;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100110 : begin
                   	state <= 10'b0011100111;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1C;
                   	IPMAdd_Z__addr_r <= 5'h11;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h10;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   end
                   10'b0011100111 : begin
                   	state <= 10'b0011101000;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h19;
                   	IPMAdd_Z__addr_r <= 5'h15;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101000 : begin
                   	state <= 10'b0011101001;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h17;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z__addr_r <= 5'h15;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101001 : begin
                   	state <= 10'b0011101010;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h15;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z__addr_r <= 5'h13;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101010 : begin
                   	state <= 10'b0011101011;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h13;
                   	IPMAdd_Z__addr_r <= 5'hD;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h14;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101011 : begin
                   	state <= 10'b0011101100;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h14;
                   	IPMAdd_Z__addr_r <= 5'hC;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   end
                   10'b0011101100 : begin
                   	state <= 10'b0011101101;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h12;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h9;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   end
                   10'b0011101101 : begin
                   	state <= 10'b0011101110;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'h8;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101110 : begin
                   	state <= 10'b0011101111;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101111 : begin
                   	state <= 10'b0011110000;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110000 : begin
                   	state <= 10'b0011110001;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110001 : begin
                   	state <= 10'b0011110010;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110010 : begin
                   	state <= 10'b0011110011;
                   	IPMAdd_Z__addr_r <= 5'h5;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h4;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   end
                   10'b0011110011 : begin
                   	state <= 10'b0011110100;
                   	round_pt[6*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   end
                   10'b0011110100 : begin
                   	state <= 10'b0011110101;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h1E;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h1D;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110101 : begin
                   	state <= 10'b0011110110;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110110 : begin
                   	state <= 10'b0011110111;
                   	round_pt[9*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h1C;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h1B;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110111 : begin
                   	state <= 10'b0011111000;
                   	IPMAdd_Z__addr_r <= 5'h1A;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h19;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111000 : begin
                   	state <= 10'b0011111001;
                   	round_pt[12*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h18;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h17;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111001 : begin
                   	state <= 10'b0011111010;
                   	round_pt[5*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h16;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h15;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111010 : begin
                   	state <= 10'b0011111011;
                   	round_pt[15*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h14;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h13;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111011 : begin
                   	state <= 10'b0011111100;
                   	round_pt[16*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h12;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h11;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111100 : begin
                   	state <= 10'b0011111101;
                   	round_pt[8*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111101 : begin
                   	state <= 10'b0011111110;
                   	round_pt[7*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'hE;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'hD;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111110 : begin
                   	state <= 10'b0011111111;
                   	round_pt[11*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'hC;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111111 : begin
                   	state <= 10'b0100000000;
                   	round_pt[2*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h9;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0100000000 : begin
                   	state <= 10'b0100000001;
                   	round_pt[3*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h8;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0100000001 : begin
                   	state <= 10'b0100000010;
                   	round_pt[10*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0100000010 : begin
                   	state <= 10'b0100000011;
                   	round_pt[14*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0100000011 : begin
                   	state <= 10'b0100000100;
                   	round_pt[13*8*v-1 -: 8*v] <= IPMAdd_P;
                   	round_count <= round_count + 1; // sen_ding this two cycles early to receive values from ks earlier
                   	IPMAdd_Z__addr_r <= 5'h2;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_add;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0100000100 : begin
                   	state <= 10'b0100000101;
                   	round_pt[1*8*v-1 -: 8*v] <= IPMAdd_P;
                   end
                   10'b0100000101 : begin
                   	state <= {is_last, 9'b000000000};
                   	round_pt[4*8*v-1 -: 8*v] <= IPMAdd_P;
                   end
                   // LAST ROUND STARTS HERE
                   10'b1000000000 : begin
                   	state <= 10'b1000000001;
                   	IPMAdd_Z_addr_r <= 5'h10; // addr of byte F
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h10; // addr of byte F
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   end
                   10'b1000000001 : begin
                   	state <= 10'b1000000010;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hF; // addr of byte E
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hF; // addr of byte E
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000000010 : begin
                   	state <= 10'b1000000011;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hE; // addr of byte D
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hE; // addr of byte D
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h5;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000000011 : begin
                   	state <= 10'b1000000100;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hD; // addr of byte C
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hD; // addr of byte C
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMMult_addr_w <= 5'h15;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h8;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h15;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000000100 : begin
                   	state <= 10'b1000000101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hC; // addr of byte B
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hC; // addr of byte B
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h4;
                   	IPMMult_addr_w <= 5'h19;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h5;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000000101 : begin
                   	state <= 10'b1000000110;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hB; // addr of byte A
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hB; // addr of byte A
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMMult_addr_w <= 5'h16;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h10;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000000110 : begin
                   	state <= 10'b1000000111;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'hA; // addr of byte 9
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'hA; // addr of byte 9
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h6;
                   	IPMMult_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h15;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h19;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000000111 : begin
                   	state <= 10'b1000001000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h9; // addr of byte 8
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h9; // addr of byte 8
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMult_addr_w <= 5'h15;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h8;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000001000 : begin
                   	state <= 10'b1000001001;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h8; // addr of byte 7
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h8; // addr of byte 7
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMult_addr_w <= 5'h13;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h4;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000001001 : begin
                   	state <= 10'b1000001010;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h7; // addr of byte 6
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h7; // addr of byte 6
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h9;
                   	IPMMult_addr_w <= 5'h9;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h5;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000001010 : begin
                   	state <= 10'b1000001011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h6; // addr of byte 5
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h6; // addr of byte 5
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMult_addr_w <= 5'h1C;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h10;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000001011 : begin
                   	state <= 10'b1000001100;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h5; // addr of byte 4
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h5; // addr of byte 4
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMMult_addr_w <= 5'hE;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMMult_Z_addr_r <= 5'h3;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h6;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h15;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000001100 : begin
                   	state <= 10'b1000001101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h4; // addr of byte 3
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h4; // addr of byte 3
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMult_addr_w <= 5'h15;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000001101 : begin
                   	state <= 10'b1000001110;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h3; // addr of byte 2
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h3; // addr of byte 2
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hC;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h19;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000001110 : begin
                   	state <= 10'b1000001111;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h2; // addr of byte 1
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h2; // addr of byte 1
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hD;
                   	IPMMult_addr_w <= 5'h19;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h7;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000001111 : begin
                   	state <= 10'b1000010000;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z_addr_r <= 5'h1; // addr of byte 0
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	IPMAdd_Z__addr_r <= 5'h1; // addr of byte 0
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMult_addr_w <= 5'h12;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h8;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000010000 : begin
                   	state <= 10'b1000010001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMult_addr_w <= 5'h18;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h4;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000010001 : begin
                   	state <= 10'b1000010010;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h9;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000010010 : begin
                   	state <= 10'b1000010011;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h17;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h8;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h1C;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000010011 : begin
                   	state <= 10'b1000010100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h5;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000010100 : begin
                   	state <= 10'b1000010101;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hC;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hA;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000010101 : begin
                   	state <= 10'b1000010110;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h1B;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h10;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000010110 : begin
                   	state <= 10'b1000010111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h1A;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMSquare_Z_addr_r <= 5'h15;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000010111 : begin
                   	state <= 10'b1000011000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h6;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000011000 : begin
                   	state <= 10'b1000011001;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMMult_Z_addr_r <= 5'hA;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hB;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000011001 : begin
                   	state <= 10'b1000011010;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h14;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMMult_Z_addr_r <= 5'hA;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hC;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h19;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000011010 : begin
                   	state <= 10'b1000011011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h19;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000011011 : begin
                   	state <= 10'b1000011100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hD;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h12;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000011100 : begin
                   	state <= 10'b1000011101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h11;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h7;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000011101 : begin
                   	state <= 10'b1000011110;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hE;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000011110 : begin
                   	state <= 10'b1000011111;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hD;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h9;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h18;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000011111 : begin
                   	state <= 10'b1000100000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h9;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h8;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000100000 : begin
                   	state <= 10'b1000100001;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h2;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hF;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h17;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000100001 : begin
                   	state <= 10'b1000100010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hF;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h9;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000100010 : begin
                   	state <= 10'b1000100011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000100011 : begin
                   	state <= 10'b1000100100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1C;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h1B;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000100100 : begin
                   	state <= 10'b1000100101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h1C;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hA;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000100101 : begin
                   	state <= 10'b1000100110;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMMult_Z_addr_r <= 5'h3;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h16;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h1A;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000100110 : begin
                   	state <= 10'b1000100111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h16;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMMult_Z_addr_r <= 5'h3;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h10;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h16;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000100111 : begin
                   	state <= 10'b1000101000;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	can_supply_last <= 1'b1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMult_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h15;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h14;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000101000 : begin
                   	state <= 10'b1000101001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMMult_addr_w <= 5'h15;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hB;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000101001 : begin
                   	state <= 10'b1000101010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h5;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMSquare_Z_addr_r <= 5'h19;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000101010 : begin
                   	state <= 10'b1000101011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMMult_Z_addr_r <= 5'hD;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hC;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000101011 : begin
                   	state <= 10'b1000101100;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h12;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h11;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000101100 : begin
                   	state <= 10'b1000101101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h12;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hD;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000101101 : begin
                   	state <= 10'b1000101110;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMMult_Z_addr_r <= 5'h4;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hE;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000101110 : begin
                   	state <= 10'b1000101111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h9;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000101111 : begin
                   	state <= 10'b1000110000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h18;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000110000 : begin
                   	state <= 10'b1000110001;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h18;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h17;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000110001 : begin
                   	state <= 10'b1000110010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h17;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hF;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000110010 : begin
                   	state <= 10'b1000110011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMSquare_Z_addr_r <= 5'h1C;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000110011 : begin
                   	state <= 10'b1000110100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000110100 : begin
                   	state <= 10'b1000110101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMult_Z_addr_r <= 5'h10;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1B;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h16;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000110101 : begin
                   	state <= 10'b1000110110;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h16;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000110110 : begin
                   	state <= 10'b1000110111;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h10;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'h3;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1A;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h15;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000110111 : begin
                   	state <= 10'b1000111000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMMult_addr_w <= 5'h15;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111000 : begin
                   	state <= 10'b1000111001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMult_Z_addr_r <= 5'hF;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h14;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111001 : begin
                   	state <= 10'b1000111010;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h14;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMMult_Z_addr_r <= 5'hA;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h13;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111010 : begin
                   	state <= 10'b1000111011;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h13;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMMult_Z_addr_r <= 5'hD;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h19;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h13;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h12;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000111011 : begin
                   	state <= 10'b1000111100;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMult_addr_w <= 5'h12;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111100 : begin
                   	state <= 10'b1000111101;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h11;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111101 : begin
                   	state <= 10'b1000111110;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h11;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMMult_Z_addr_r <= 5'h4;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hD;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111110 : begin
                   	state <= 10'b1000111111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hD;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMSquare_Z_addr_r <= 5'h18;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000111111 : begin
                   	state <= 10'b1001000000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMSquare_Z_addr_r <= 5'h17;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001000000 : begin
                   	state <= 10'b1001000001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001000001 : begin
                   	state <= 10'b1001000010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hF;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001000010 : begin
                   	state <= 10'b1001000011;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hF;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMMult_Z_addr_r <= 5'hB;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hE;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001000011 : begin
                   	state <= 10'b1001000100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hE;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001000100 : begin
                   	state <= 10'b1001000101;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h16;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001000101 : begin
                   	state <= 10'b1001000110;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h10;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001000110 : begin
                   	state <= 10'b1001000111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMSquare_Z_addr_r <= 5'h15;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001000111 : begin
                   	state <= 10'b1001001000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMSquare_Z_addr_r <= 5'h14;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001001000 : begin
                   	state <= 10'b1001001001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMSquare_Z_addr_r <= 5'h13;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001001001 : begin
                   	state <= 10'b1001001010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001001010 : begin
                   	state <= 10'b1001001011;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h12;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001001011 : begin
                   	state <= 10'b1001001100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMSquare_Z_addr_r <= 5'h11;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001001100 : begin
                   	state <= 10'b1001001101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001001101 : begin
                   	state <= 10'b1001001110;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMMult_Z_addr_r <= 5'h9;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h10;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001001110 : begin
                   	state <= 10'b1001001111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'hD;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001001111 : begin
                   	state <= 10'b1001010000;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010000 : begin
                   	state <= 10'b1001010001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hD;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001010001 : begin
                   	state <= 10'b1001010010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001010010 : begin
                   	state <= 10'b1001010011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010011 : begin
                   	state <= 10'b1001010100;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'h2;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hC;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010100 : begin
                   	state <= 10'b1001010101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMult_addr_w <= 5'hC;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010101 : begin
                   	state <= 10'b1001010110;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h10;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010110 : begin
                   	state <= 10'b1001010111;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMult_Z_addr_r <= 5'h3;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h7;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010111 : begin
                   	state <= 10'b1001011000;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hC;
                   	IPMMult_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011000 : begin
                   	state <= 10'b1001011001;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011001 : begin
                   	state <= 10'b1001011010;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011010 : begin
                   	state <= 10'b1001011011;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'hD;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hA;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011011 : begin
                   	state <= 10'b1001011100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMult_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011100 : begin
                   	state <= 10'b1001011101;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001011101 : begin
                   	state <= 10'b1001011110;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011110 : begin
                   	state <= 10'b1001011111;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hD;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011111 : begin
                   	state <= 10'b1001100000;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hD;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMMult_Z_addr_r <= 5'h4;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h2;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100000 : begin
                   	state <= 10'b1001100001;
                   	IPMMult_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_addr_w <= 5'h2;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMMult_Z_addr_r <= 5'hC;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h8;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100001 : begin
                   	state <= 10'b1001100010;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMMult_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100010 : begin
                   	state <= 10'b1001100011;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'h9;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100011 : begin
                   	state <= 10'b1001100100;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001100100 : begin
                   	state <= 10'b1001100101;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h10;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100101 : begin
                   	state <= 10'b1001100110;
                   	IPMMultConst_const <= 8'h5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hC;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'hB;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'hB;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001100110 : begin
                   	state <= 10'b1001100111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hC;
                   	IPMMult_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100111 : begin
                   	state <= 10'b1001101000;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'h5;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h6;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101000 : begin
                   	state <= 10'b1001101001;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMult_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMult_Z_addr_r <= 5'hA;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h5;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101001 : begin
                   	state <= 10'b1001101010;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMult_addr_w <= 5'h5;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001101010 : begin
                   	state <= 10'b1001101011;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101011 : begin
                   	state <= 10'b1001101100;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMult_Z_addr_r <= 5'h6;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h4;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101100 : begin
                   	state <= 10'b1001101101;
                   	IPMMultConst_const <= 8'h5;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMMult_addr_w <= 5'h4;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'h8;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h3;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101101 : begin
                   	state <= 10'b1001101110;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMult_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101110 : begin
                   	state <= 10'b1001101111;
                   	IPMMultConst_const <= 8'h9;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h4;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hD;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMult_Z_addr_r <= 5'h9;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h9;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001101111 : begin
                   	state <= 10'b1001110000;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'hD;
                   	IPMMult_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001110000 : begin
                   	state <= 10'b1001110001;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h9;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001110001 : begin
                   	state <= 10'b1001110010;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'h9;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMult_Z_addr_r <= 5'h7;
                   	IPMMult_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMMult_Z__addr_r <= 5'h1;
                   	IPMMult_Z__addr_r_BRAM <= BRAM_mul;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001110010 : begin
                   	state <= 10'b1001110011;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMult_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMult_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001110011 : begin
                   	state <= 10'b1001110100;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001110100 : begin
                   	state <= 10'b1001110101;
                   	IPMMultConst_const <= 8'h8f;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mask; // take from IPMMask
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_mc;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001110101 : begin
                   	state <= 10'b1001110110;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h10;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001110110 : begin
                   	state <= 10'b1001110111;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hC;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001110111 : begin
                   	state <= 10'b1001111000;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hC;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001111000 : begin
                   	state <= 10'b1001111001;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001111001 : begin
                   	state <= 10'b1001111010;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001111010 : begin
                   	state <= 10'b1001111011;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001111011 : begin
                   	state <= 10'b1001111100;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001111100 : begin
                   	state <= 10'b1001111101;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001111101 : begin
                   	state <= 10'b1001111110;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h4;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001111110 : begin
                   	state <= 10'b1001111111;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h4;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hD;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001111111 : begin
                   	state <= 10'b1010000000;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hD;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000000 : begin
                   	state <= 10'b1010000001;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h9;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000001 : begin
                   	state <= 10'b1010000010;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h9;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1010000010 : begin
                   	state <= 10'b1010000011;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000011 : begin
                   	state <= 10'b1010000100;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'h10;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h10;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000100 : begin
                   	state <= 10'b1010000101;
                   	IPMMultConst_const <= 8'h5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000101 : begin
                   	state <= 10'b1010000110;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000110 : begin
                   	state <= 10'b1010000111;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hC;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000111 : begin
                   	state <= 10'b1010001000;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hC;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001000 : begin
                   	state <= 10'b1010001001;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001001 : begin
                   	state <= 10'b1010001010;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001010 : begin
                   	state <= 10'b1010001011;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001011 : begin
                   	state <= 10'b1010001100;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001100 : begin
                   	state <= 10'b1010001101;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001101 : begin
                   	state <= 10'b1010001110;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h4;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001110 : begin
                   	state <= 10'b1010001111;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h4;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hD;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001111 : begin
                   	state <= 10'b1010010000;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hD;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010000 : begin
                   	state <= 10'b1010010001;
                   	IPMMultConst_const <= 8'h9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h9;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010001 : begin
                   	state <= 10'b1010010010;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h9;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010010 : begin
                   	state <= 10'b1010010011;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h10;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010011 : begin
                   	state <= 10'b1010010100;
                   	IPMMultConst_const <= 8'h9;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h10;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h10;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010100 : begin
                   	state <= 10'b1010010101;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010101 : begin
                   	state <= 10'b1010010110;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h10;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010110 : begin
                   	state <= 10'b1010010111;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h10;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hC;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010111 : begin
                   	state <= 10'b1010011000;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r <= 5'h4; // addr of byte 3
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hC;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z_addr_r <= 5'h10;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011000 : begin
                   	state <= 10'b1010011001;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011001 : begin
                   	state <= 10'b1010011010;
                   	round_pt[4*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011010 : begin
                   	state <= 10'b1010011011;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'hF;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011011 : begin
                   	state <= 10'b1010011100;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011100 : begin
                   	state <= 10'b1010011101;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011101 : begin
                   	state <= 10'b1010011110;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011110 : begin
                   	state <= 10'b1010011111;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h4;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011111 : begin
                   	state <= 10'b1010100000;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h4;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hD;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100000 : begin
                   	state <= 10'b1010100001;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hD;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100001 : begin
                   	state <= 10'b1010100010;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h9;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100010 : begin
                   	state <= 10'b1010100011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h9;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100011 : begin
                   	state <= 10'b1010100100;
                   	IPMMultConst_const <= 8'hf9;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'hE;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100100 : begin
                   	state <= 10'b1010100101;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100101 : begin
                   	state <= 10'b1010100110;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100110 : begin
                   	state <= 10'b1010100111;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hC;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hF;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100111 : begin
                   	state <= 10'b1010101000;
                   	IPMMultConst_const <= 8'h25;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hC;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'hF;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hF;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101000 : begin
                   	state <= 10'b1010101001;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101001 : begin
                   	state <= 10'b1010101010;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101010 : begin
                   	state <= 10'b1010101011;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101011 : begin
                   	state <= 10'b1010101100;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hF;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101100 : begin
                   	state <= 10'b1010101101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101101 : begin
                   	state <= 10'b1010101110;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r <= 5'h7; // addr of byte 6
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z_addr_r <= 5'hF;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101110 : begin
                   	state <= 10'b1010101111;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'hD;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'hD;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101111 : begin
                   	state <= 10'b1010110000;
                   	round_pt[7*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hD;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h4;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hE;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110000 : begin
                   	state <= 10'b1010110001;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h4;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'hE;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hE;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110001 : begin
                   	state <= 10'b1010110010;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h9;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110010 : begin
                   	state <= 10'b1010110011;
                   	IPMMultConst_const <= 8'h25;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h9;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110011 : begin
                   	state <= 10'b1010110100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110100 : begin
                   	state <= 10'b1010110101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110101 : begin
                   	state <= 10'b1010110110;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hE;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'hC;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'hC;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110110 : begin
                   	state <= 10'b1010110111;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hC;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110111 : begin
                   	state <= 10'b1010111000;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'hB;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111000 : begin
                   	state <= 10'b1010111001;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r <= 5'hA; // addr of byte 9
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z_addr_r <= 5'hE;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hD;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111001 : begin
                   	state <= 10'b1010111010;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'hD;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hD;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111010 : begin
                   	state <= 10'b1010111011;
                   	round_pt[10*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111011 : begin
                   	state <= 10'b1010111100;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h6;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'hA;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111100 : begin
                   	state <= 10'b1010111101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111101 : begin
                   	state <= 10'b1010111110;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h4;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111110 : begin
                   	state <= 10'b1010111111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hD;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h1;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hC;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111111 : begin
                   	state <= 10'b1011000000;
                   	IPMMultConst_const <= 8'hf4;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hD;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'hC;
                   	IPMAdd_Z__addr_r <= 5'h9;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h9;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hC;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'hB;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000000 : begin
                   	state <= 10'b1011000001;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h9;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'hB;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hB;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000001 : begin
                   	state <= 10'b1011000010;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'h8;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000010 : begin
                   	state <= 10'b1011000011;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000011 : begin
                   	state <= 10'b1011000100;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r <= 5'hD; // addr of byte C
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z_addr_r <= 5'hD;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'hA;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000100 : begin
                   	state <= 10'b1011000101;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMSquare_addr_w <= 5'hA;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'hA;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000101 : begin
                   	state <= 10'b1011000110;
                   	round_pt[13*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hC;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000110 : begin
                   	state <= 10'b1011000111;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hC;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h9;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000111 : begin
                   	state <= 10'b1011001000;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hB;
                   	IPMSquare_addr_w <= 5'h9;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h9;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001000 : begin
                   	state <= 10'b1011001001;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h8;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001001 : begin
                   	state <= 10'b1011001010;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h8;
                   	IPMAdd_Z__addr_r <= 5'h5;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h8;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001010 : begin
                   	state <= 10'b1011001011;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMSquare_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMSquare_Z_addr_r <= 5'h7;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001011 : begin
                   	state <= 10'b1011001100;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'hA;
                   	IPMSquare_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h4;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h7;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h6;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001100 : begin
                   	state <= 10'b1011001101;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r <= 5'h10; // addr of byte F
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h4;
                   	IPMMultConst_addr_w <= 5'h7;
                   	IPMSquare_addr_w <= 5'h6;
                   	IPMAdd_Z_addr_r <= 5'hC;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h6;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h5;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001101 : begin
                   	state <= 10'b1011001110;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h6;
                   	IPMSquare_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h5;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h4;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001110 : begin
                   	state <= 10'b1011001111;
                   	round_pt[16*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r <= 5'h3; // addr of byte 2
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMMultConst_addr_w <= 5'h5;
                   	IPMSquare_addr_w <= 5'h4;
                   	IPMAdd_Z_addr_r <= 5'hB;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h4;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h3;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001111 : begin
                   	state <= 10'b1011010000;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMMultConst_addr_w <= 5'h4;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h9;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h2;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011010000 : begin
                   	state <= 10'b1011010001;
                   	round_pt[3*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h9;
                   	IPMMultConst_addr_w <= 5'h3;
                   	IPMSquare_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h2;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h3;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	IPMSquare_Z_addr_r <= 5'h1;
                   	IPMSquare_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011010001 : begin
                   	state <= 10'b1011010010;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMSquare_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMMultConst_addr_w <= 5'h2;
                   	IPMSquare_addr_w <= 5'h2;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   	IPMMultConst_Z_addr_r <= 5'h2;
                   	IPMMultConst_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011010010 : begin
                   	state <= 10'b1011010011;
                   	IPMMultConst_const <= 8'hb5;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMMultConst_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h8;
                   	IPMMultConst_addr_w <= 5'h1;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_sq;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011010011 : begin
                   	state <= 10'b1011010100;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r <= 5'h6; // addr of byte 5
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMAdd_Z_addr_r <= 5'hA;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011010100 : begin
                   	state <= 10'b1011010101;
                   	IPMAdd_Z__addr_r <= 5'h7;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011010101 : begin
                   	state <= 10'b1011010110;
                   	round_pt[6*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h7;
                   	IPMAdd_Z__addr_r <= 5'h6;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011010110 : begin
                   	state <= 10'b1011010111;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h6;
                   	IPMAdd_Z__addr_r <= 5'h5;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011010111 : begin
                   	state <= 10'b1011011000;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h5;
                   	IPMAdd_Z__addr_r <= 5'h4;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h4;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011000 : begin
                   	state <= 10'b1011011001;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r <= 5'h9; // addr of byte 8
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h4;
                   	IPMAdd_Z_addr_r <= 5'h9;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011001 : begin
                   	state <= 10'b1011011010;
                   	IPMAdd_Z__addr_r <= 5'h3;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011010 : begin
                   	state <= 10'b1011011011;
                   	round_pt[9*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_addr_w <= 5'h3;
                   	IPMAdd_Z__addr_r <= 5'h2;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011011 : begin
                   	state <= 10'b1011011100;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r <= 5'hC; // addr of byte B
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h2;
                   	IPMAdd_Z_addr_r <= 5'h8;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011100 : begin
                   	state <= 10'b1011011101;
                   	IPMAdd_Z__addr_r <= 5'h1;
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_mc;
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011101 : begin
                   	state <= 10'b1011011110;
                   	round_pt[12*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_BRAM_en <= 1;
                   	IPMAdd_Z__addr_r <= 5'hF; // addr of byte E
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_addr_w <= 5'h1;
                   	IPMAdd_Z_addr_r <= 5'h7;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011110 : begin
                   	state <= 10'b1011011111;
                   	IPMAdd_Z__addr_r <= 5'h2; // addr of byte 1
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_Z_addr_r <= 5'h6;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011111 : begin
                   	state <= 10'b1011100000;
                   	round_pt[15*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h5; // addr of byte 4
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_Z_addr_r <= 5'h5;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011100000 : begin
                   	state <= 10'b1011100001;
                   	round_pt[2*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h8; // addr of byte 7
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_Z_addr_r <= 5'h4;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011100001 : begin
                   	state <= 10'b1011100010;
                   	round_pt[5*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'hB; // addr of byte A
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_Z_addr_r <= 5'h3;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011100010 : begin
                   	state <= 10'b1011100011;
                   	round_pt[8*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'hE; // addr of byte D
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_Z_addr_r <= 5'h2;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011100011 : begin
                   	state <= 10'b1011100100;
                   	round_pt[11*8*v-1 -: 8*v] <= IPMAdd_P;
                   	IPMAdd_Z__addr_r <= 5'h1; // addr of byte 0
                   	IPMAdd_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	IPMAdd_Z_addr_r <= 5'h1;
                   	IPMAdd_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011100100 : begin
                   	state <= 10'b1011100101;
                   	round_pt[14*8*v-1 -: 8*v] <= IPMAdd_P;
                   end
                   10'b1011100101 : begin
                   	state <= 10'b1111111100;
                   	round_pt[1*8*v-1 -: 8*v] <= IPMAdd_P;
                   	is_busy <= 1'b0;
                   end
                   default : begin
                   	state <= 10'b1111111100;
                   end
                endcase
            end
        end
    end


endmodule