/**
 * Module: identity8
 * 
 * TODO: Add module documentation
 */
module identity8 (
	input	[7:0]	x,
	output	[7:0]	y
);
	
	assign x = y;


endmodule


