/****************************************************************************

 * roundAES.v

 ****************************************************************************/



/**

 * Module: roundAES

 * 

 * TODO: Add module documentation

 */
module roundAES (
	input  clk,
	input  rst,
	input  en,
	input [16*8-1:0] plaintext,
	input [16*8-1:0] round_ks,
	output reg can_supply_last,
	output [3:0] current_round,
	output [16*8-1:0] ciphertext,
	output reg is_busy
);

    // just have this so you do not need to replace all the "v*" and "*v"
    parameter v = 1;
    // bram adresses
    parameter BRAM_mul = 3'b000;
    parameter BRAM_add = 3'b001;
    parameter BRAM_sq = 3'b010;
    parameter BRAM_mc = 3'b011;
    parameter BRAM_PT = 3'b100;
    parameter BRAM_KS = 3'b101;
    parameter BRAM_mask = 3'b110;
    parameter BRAM_DEFAULT = 3'b111;


	wire RNGisReady = 1;
	reg RNGenable;
	reg RNGreseed;
	reg RNGisInit = 0;


    reg [16*8-1:0] round_pt;

	//==============================
	// wires :
	//==============================


	wire  [8-1:0] Square_Z;
	wire [8-1:0] Square_P;
	wire  [8-1:0] Mult_Z;
	wire  [8-1:0] Mult_Z_;
	wire [8-1:0] Mult_P;
	wire  [8-1:0] Add_Z;
	wire  [8-1:0] Add_Z_;
	wire [8-1:0] Add_P;
	wire [8-1:0] Mask_R;
	wire  [8-1:0] MultConst_Z;
	reg  [8-1:0] MultConst_const;
	wire [8-1:0] MultConst_P;


	reg  [10-1:0] state;
	reg  [3:0] round_count;
	assign current_round = round_count;

	//==============================
	// IO :
	//==============================
	assign ciphertext = round_pt;

	//==============================
	// modules :
	//==============================
	square8 square8(
		.a(Square_Z),
		.b(Square_P)
	);

	gmul8 gmul8(
		.x(Mult_Z),
		.y(Mult_Z_),
		.xy(Mult_P)
	);

	gadd8 gadd8(
		.x(Add_Z),
		.y(Add_Z_),
		.xy(Add_P)
	);

	identity8 identity8(
		.x(8'h63),
		.y(Mask_R)
	);

    // multConst is done by a normal gmul8 module
	gmul8 gmul8_mc(
		.x(MultConst_Z),
		.y(MultConst_const),
		.xy(MultConst_P)
	);



	reg Add_BRAM_en;
	reg Mult_BRAM_en;
	reg MultConst_BRAM_en;
	reg Square_BRAM_en;
	reg [4:0] Add_addr_w;
	reg [4:0] Mult_addr_w;
	reg [4:0] MultConst_addr_w;
	reg [4:0] Square_addr_w;

    reg [4:0] Add_Z_addr_r;
    reg [4:0] Add_Z__addr_r;
    reg [4:0] Mult_Z_addr_r;
    reg [4:0] Mult_Z__addr_r;
    reg [4:0] MultConst_Z_addr_r;
    reg [4:0] Square_Z_addr_r;

    reg [2:0] Add_Z_addr_r_BRAM;
    reg [2:0] Add_Z__addr_r_BRAM;
    reg [2:0] Mult_Z_addr_r_BRAM;
    reg [2:0] Mult_Z__addr_r_BRAM;
    reg [2:0] MultConst_Z_addr_r_BRAM;
    reg [2:0] Square_Z_addr_r_BRAM;

    Bank #(.addr_bits(5), .debug(1)) Bank (
         .DEBUG_STATE(state),
         .clk(clk),
         .en(en),
         .plaintext(round_pt),
         .round_ks(round_ks),
         .add_en(Add_BRAM_en),
         .mul_en(Mult_BRAM_en),
         .mc_en(MultConst_BRAM_en),
         .sq_en(Square_BRAM_en),
         .add_addr_w(Add_addr_w),
         .mul_addr_w(Mult_addr_w),
         .mc_addr_w(MultConst_addr_w),
         .sq_addr_w(Square_addr_w),
         .add_val_w(Add_P),
         .mul_val_w(Mult_P),
         .mc_val_w(MultConst_P),
         .sq_val_w(Square_P),
         .mask_val_w(Mask_R),
         .add0_addr_r(Add_Z_addr_r),
         .add1_addr_r(Add_Z__addr_r),
         .mul0_addr_r(Mult_Z_addr_r),
         .mul1_addr_r(Mult_Z__addr_r),
         .mc_addr_r(MultConst_Z_addr_r),
         .sq_addr_r(Square_Z_addr_r),
         .add0_r_BRAM(Add_Z_addr_r_BRAM),
         .add1_r_BRAM(Add_Z__addr_r_BRAM),
         .mul0_r_BRAM(Mult_Z_addr_r_BRAM),
         .mul1_r_BRAM(Mult_Z__addr_r_BRAM),
         .mc_r_BRAM(MultConst_Z_addr_r_BRAM),
         .sq_r_BRAM(Square_Z_addr_r_BRAM),
         .add0_out(Add_Z),
         .add1_out(Add_Z_),
         .mul0_out(Mult_Z),
         .mul1_out(Mult_Z_),
         .mc_out(MultConst_Z),
         .sq_out(Square_Z)
    );




	//==============================
	// control :
	//==============================


	wire is_last = (round_count == 10);
	always @(posedge clk) begin
		if (!rst) begin
			state <= 10'b1111111111;
			is_busy <= 1;
		end
		else begin
            if(!en) begin
                state <= 10'b1111111111;
					 is_busy <= 1;
            end else begin


                // these are important!!!
                Add_BRAM_en <= 0;
                Mult_BRAM_en <= 0;
                MultConst_BRAM_en <= 0;
                Square_BRAM_en <= 0;
                Add_Z_addr_r_BRAM <= BRAM_DEFAULT;
                Add_Z__addr_r_BRAM <= BRAM_DEFAULT;
                Mult_Z_addr_r_BRAM <= BRAM_DEFAULT;
                Mult_Z__addr_r_BRAM <= BRAM_DEFAULT;
                Square_Z_addr_r_BRAM <= BRAM_DEFAULT;
                MultConst_Z_addr_r_BRAM <= BRAM_DEFAULT;
                MultConst_const <= 8'h0;
                // 0 address is not in use
                Square_addr_w <= 8'h0;
                Mult_addr_w <= 8'h0;
                Add_addr_w <= 8'h0;
                MultConst_addr_w <= 8'h0;

                // FSM
                case(state)                    // reset RNG
                    10'b1111111111 : begin
                        can_supply_last <= 0;
                        RNGreseed <= 1;
                        RNGenable <= 1;
                        state <= 10'b1111111110;
                        round_count <= 1;
                        round_pt <= plaintext[1*16*v*8-1:0*16*v*8];
                        is_busy <= 1;
                    end
                    // wait until RNG is ready
                    10'b1111111110 : begin
                        RNGreseed <= 0;
                        if (RNGisReady) begin
                            state <= 10'b0000000000;
                        end else begin
                            state <= 10'b1111111110;
                        end
                    end
                    // rounds 1-9 start here
                   10'b0000000000 : begin
                   	state <= 10'b0000000001;
                   	Add_Z_addr_r <= 5'h10; // addr of byte F
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h10; // addr of byte F
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   end
                   10'b0000000001 : begin
                   	state <= 10'b0000000010;
                   	Add_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hF; // addr of byte E
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hF; // addr of byte E
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h11;
                   	Square_Z_addr_r <= 5'h11;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000000010 : begin
						 
                   	state <= 10'b0000000011;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hE; // addr of byte D
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hE; // addr of byte D
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h11;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000000011 : begin
						 
                   	
                   	state <= 10'b0000000100;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hD; // addr of byte C
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hD; // addr of byte C
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hE;
                   	Mult_addr_w <= 5'h15;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hA;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h15;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000000100 : begin
						 
                   	
                   	state <= 10'b0000000101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hC; // addr of byte B
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hC; // addr of byte B
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h3;
                   	Mult_addr_w <= 5'h19;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h11;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000000101 : begin
						 
                   	
                   	state <= 10'b0000000110;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hB; // addr of byte A
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hB; // addr of byte A
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h11;
                   	Mult_addr_w <= 5'h16;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hE;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000000110 : begin
						 
                   	
                   	
                   	state <= 10'b0000000111;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hA; // addr of byte 9
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hA; // addr of byte 9
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h1;
                   	Mult_addr_w <= 5'h8;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h15;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h19;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000000111 : begin
						 
                   	
                   	
                   	state <= 10'b0000001000;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h9; // addr of byte 8
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h9; // addr of byte 8
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h16;
                   	Mult_addr_w <= 5'h15;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hA;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000001000 : begin
						 
                   	
                   	
                   	state <= 10'b0000001001;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h8; // addr of byte 7
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h8; // addr of byte 7
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hA;
                   	Mult_addr_w <= 5'h13;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h3;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h11;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000001001 : begin
						 
                   	
                   	
                   	state <= 10'b0000001010;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h7; // addr of byte 6
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h7; // addr of byte 6
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hF;
                   	Mult_addr_w <= 5'h9;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h11;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000001010 : begin
						 
                   	
                   	
                   	state <= 10'b0000001011;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h6; // addr of byte 5
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h6; // addr of byte 5
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h13;
                   	Mult_addr_w <= 5'h1C;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hE;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000001011 : begin
						 
                   	
                   	
                   	state <= 10'b0000001100;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h5; // addr of byte 4
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h5; // addr of byte 4
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hE;
                   	Mult_addr_w <= 5'hE;
                   	Square_addr_w <= 5'h3;
                   	Mult_Z_addr_r <= 5'h3;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h15;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000001100 : begin
						 
                   	
                   	
                   	state <= 10'b0000001101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h4; // addr of byte 3
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h4; // addr of byte 3
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h2;
                   	Mult_addr_w <= 5'h15;
                   	Square_addr_w <= 5'h3;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000001101 : begin
						 
                   	
                   	
                   	state <= 10'b0000001110;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h3; // addr of byte 2
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h3; // addr of byte 2
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h8;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h19;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h16;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000001110 : begin
						 
                   	
                   	
                   	state <= 10'b0000001111;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h2; // addr of byte 1
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h2; // addr of byte 1
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h7;
                   	Mult_addr_w <= 5'h19;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h16;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000001111 : begin
						 
                   	
                   	
                   	state <= 10'b0000010000;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h1; // addr of byte 0
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h1; // addr of byte 0
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h1B;
                   	Mult_addr_w <= 5'h12;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hA;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000010000 : begin
						 
                   	
                   	
                   	state <= 10'b0000010001;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h14;
                   	Mult_addr_w <= 5'h18;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h3;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000010001 : begin
						 
                   	
                   	
                   	state <= 10'b0000010010;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h10;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hF;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000010010 : begin
                   	state <= 10'b0000010011;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h17;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h8;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h1C;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000010011 : begin
                   	state <= 10'b0000010100;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h8;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h11;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h13;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000010100 : begin
                   	state <= 10'b0000010101;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hC;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h13;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000010101 : begin
                   	state <= 10'b0000010110;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h1B;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hE;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000010110 : begin
                   	state <= 10'b0000010111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h1A;
                   	Square_addr_w <= 5'h3;
                   	Square_Z_addr_r <= 5'h15;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000010111 : begin
                   	state <= 10'b0000011000;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000011000 : begin
                   	state <= 10'b0000011001;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h7;
                   	Square_addr_w <= 5'hA;
                   	Mult_Z_addr_r <= 5'hA;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h2;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000011001 : begin
                   	state <= 10'b0000011010;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h14;
                   	Square_addr_w <= 5'hA;
                   	Mult_Z_addr_r <= 5'hA;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h8;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h19;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000011010 : begin
                   	state <= 10'b0000011011;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h19;
                   	Square_addr_w <= 5'hA;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000011011 : begin
                   	state <= 10'b0000011100;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h7;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h12;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000011100 : begin
                   	state <= 10'b0000011101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h11;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h16;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h1B;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000011101 : begin
                   	state <= 10'b0000011110;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1B;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000011110 : begin
                   	state <= 10'b0000011111;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hD;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h9;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h18;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000011111 : begin
                   	state <= 10'b0000100000;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h9;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hA;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h14;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0000100000 : begin
                   	state <= 10'b0000100001;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h2;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h14;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h17;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000100001 : begin
                   	state <= 10'b0000100010;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hF;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hF;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000100010 : begin
                   	state <= 10'b0000100011;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h8;
                   	Square_addr_w <= 5'hB;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000100011 : begin
                   	state <= 10'b0000100100;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1C;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h1B;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000100100 : begin
                   	state <= 10'b0000100101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h1C;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h13;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000100101 : begin
                   	state <= 10'b0000100110;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hB;
                   	Square_addr_w <= 5'h3;
                   	Mult_Z_addr_r <= 5'h3;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h16;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h1A;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000100110 : begin
                   	state <= 10'b0000100111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h16;
                   	Square_addr_w <= 5'h3;
                   	Mult_Z_addr_r <= 5'h3;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hE;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h16;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000100111 : begin
                   	state <= 10'b0000101000;
                   	MultConst_const <= 8'h8f;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Mult_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hF;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h15;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h14;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000101000 : begin
                   	state <= 10'b0000101001;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	Mult_addr_w <= 5'h15;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h2;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000101001 : begin
                   	state <= 10'b0000101010;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h5;
                   	Square_addr_w <= 5'hA;
                   	Square_Z_addr_r <= 5'h19;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000101010 : begin
                   	state <= 10'b0000101011;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hD;
                   	Mult_Z_addr_r <= 5'hD;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h8;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000101011 : begin
                   	state <= 10'b0000101100;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h12;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h11;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000101100 : begin
                   	state <= 10'b0000101101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h12;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h7;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000101101 : begin
                   	state <= 10'b0000101110;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h4;
                   	Mult_Z_addr_r <= 5'h4;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1B;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000101110 : begin
                   	state <= 10'b0000101111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h9;
                   	Square_addr_w <= 5'h9;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000101111 : begin
                   	state <= 10'b0000110000;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h18;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000110000 : begin
                   	state <= 10'b0000110001;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h18;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h17;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000110001 : begin
                   	state <= 10'b0000110010;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h17;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h14;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000110010 : begin
                   	state <= 10'b0000110011;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h1;
                   	Square_addr_w <= 5'hB;
                   	Square_Z_addr_r <= 5'h1C;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000110011 : begin
                   	state <= 10'b0000110100;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h2;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000110100 : begin
                   	state <= 10'b0000110101;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1B;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h16;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000110101 : begin
                   	state <= 10'b0000110110;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h16;
                   	Square_addr_w <= 5'h10;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000110110 : begin
                   	state <= 10'b0000110111;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'h3;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1A;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h15;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000110111 : begin
                   	state <= 10'b0000111000;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	Mult_addr_w <= 5'h15;
                   	Square_addr_w <= 5'h3;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111000 : begin
                   	state <= 10'b0000111001;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h14;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111001 : begin
                   	state <= 10'b0000111010;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h14;
                   	Square_addr_w <= 5'hA;
                   	Mult_Z_addr_r <= 5'hA;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h13;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111010 : begin
                   	state <= 10'b0000111011;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h13;
                   	Square_addr_w <= 5'hD;
                   	Mult_Z_addr_r <= 5'hD;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h19;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h13;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h12;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000111011 : begin
                   	state <= 10'b0000111100;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Mult_addr_w <= 5'h12;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hD;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111100 : begin
                   	state <= 10'b0000111101;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h14;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h11;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111101 : begin
                   	state <= 10'b0000111110;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h11;
                   	Square_addr_w <= 5'h4;
                   	Mult_Z_addr_r <= 5'h4;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hD;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0000111110 : begin
                   	state <= 10'b0000111111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hD;
                   	Square_addr_w <= 5'h9;
                   	Square_Z_addr_r <= 5'h18;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0000111111 : begin
                   	state <= 10'b0001000000;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h4;
                   	Square_Z_addr_r <= 5'h17;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001000000 : begin
                   	state <= 10'b0001000001;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hC;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001000001 : begin
                   	state <= 10'b0001000010;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hF;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001000010 : begin
                   	state <= 10'b0001000011;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hF;
                   	Square_addr_w <= 5'hB;
                   	Mult_Z_addr_r <= 5'hB;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hE;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001000011 : begin
                   	state <= 10'b0001000100;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hE;
                   	Square_addr_w <= 5'h2;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001000100 : begin
                   	state <= 10'b0001000101;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h10;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h16;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001000101 : begin
                   	state <= 10'b0001000110;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1B;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001000110 : begin
                   	state <= 10'b0001000111;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	Square_addr_w <= 5'h3;
                   	Square_Z_addr_r <= 5'h15;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001000111 : begin
                   	state <= 10'b0001001000;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h5;
                   	Square_Z_addr_r <= 5'h14;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001001000 : begin
                   	state <= 10'b0001001001;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hA;
                   	Square_Z_addr_r <= 5'h13;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001001001 : begin
                   	state <= 10'b0001001010;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hF;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001001010 : begin
                   	state <= 10'b0001001011;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h14;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h12;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001001011 : begin
                   	state <= 10'b0001001100;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h14;
                   	Square_addr_w <= 5'h6;
                   	Square_Z_addr_r <= 5'h11;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001001100 : begin
                   	state <= 10'b0001001101;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h8;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001001101 : begin
                   	state <= 10'b0001001110;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h9;
                   	Mult_Z_addr_r <= 5'h9;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h10;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001001110 : begin
                   	state <= 10'b0001001111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hD;
                   	Square_addr_w <= 5'h9;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001001111 : begin
                   	state <= 10'b0001010000;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h4;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010000 : begin
                   	state <= 10'b0001010001;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	Square_addr_w <= 5'hC;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001010001 : begin
                   	state <= 10'b0001010010;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h7;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001010010 : begin
                   	state <= 10'b0001010011;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hE;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010011 : begin
                   	state <= 10'b0001010100;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1B;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hC;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010100 : begin
                   	state <= 10'b0001010101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1B;
                   	Mult_addr_w <= 5'hC;
                   	Square_addr_w <= 5'h10;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010101 : begin
                   	state <= 10'b0001010110;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010110 : begin
                   	state <= 10'b0001010111;
                   	MultConst_const <= 8'h8f;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h3;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Mult_Z_addr_r <= 5'h3;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h7;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001010111 : begin
                   	state <= 10'b0001011000;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	Mult_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h5;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011000 : begin
                   	state <= 10'b0001011001;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hA;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011001 : begin
                   	state <= 10'b0001011010;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	Square_addr_w <= 5'hF;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011010 : begin
                   	state <= 10'b0001011011;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h14;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'hD;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hA;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011011 : begin
                   	state <= 10'b0001011100;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h14;
                   	Mult_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h6;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011100 : begin
                   	state <= 10'b0001011101;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h8;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001011101 : begin
                   	state <= 10'b0001011110;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h13;
                   	Square_addr_w <= 5'hD;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011110 : begin
                   	state <= 10'b0001011111;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001011111 : begin
                   	state <= 10'b0001100000;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h4;
                   	Mult_Z_addr_r <= 5'h4;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h2;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100000 : begin
                   	state <= 10'b0001100001;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h2;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h8;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100001 : begin
                   	state <= 10'b0001100010;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Mult_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h7;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100010 : begin
                   	state <= 10'b0001100011;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hE;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100011 : begin
                   	state <= 10'b0001100100;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1B;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001100100 : begin
                   	state <= 10'b0001100101;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1B;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100101 : begin
                   	state <= 10'b0001100110;
                   	MultConst_const <= 8'h5;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'hB;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hB;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001100110 : begin
                   	state <= 10'b0001100111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	Mult_addr_w <= 5'h7;
                   	Square_addr_w <= 5'hB;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001100111 : begin
                   	state <= 10'b0001101000;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h6;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101000 : begin
                   	state <= 10'b0001101001;
                   	MultConst_const <= 8'h8f;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'h2;
                   	Mult_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hA;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Mult_Z_addr_r <= 5'hA;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h5;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101001 : begin
                   	state <= 10'b0001101010;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'h16;
                   	Mult_addr_w <= 5'h5;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hF;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001101010 : begin
                   	state <= 10'b0001101011;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h14;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101011 : begin
                   	state <= 10'b0001101100;
                   	MultConst_const <= 8'h8f;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'h14;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h6;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Mult_Z_addr_r <= 5'h6;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h4;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101100 : begin
                   	state <= 10'b0001101101;
                   	MultConst_const <= 8'h5;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h11;
                   	Mult_addr_w <= 5'h4;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h13;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'h8;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h3;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101101 : begin
                   	state <= 10'b0001101110;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'h13;
                   	Mult_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hD;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001101110 : begin
                   	state <= 10'b0001101111;
                   	MultConst_const <= 8'h9;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'h9;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h9;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001101111 : begin
                   	state <= 10'b0001110000;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'h7;
                   	Mult_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h9;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001110000 : begin
                   	state <= 10'b0001110001;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1C;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001110001 : begin
                   	state <= 10'b0001110010;
                   	MultConst_const <= 8'h8f;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h7;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Mult_Z_addr_r <= 5'h7;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001110010 : begin
                   	state <= 10'b0001110011;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h15;
                   	Mult_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001110011 : begin
                   	state <= 10'b0001110100;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1B;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001110100 : begin
                   	state <= 10'b0001110101;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'h1B;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hC;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001110101 : begin
                   	state <= 10'b0001110110;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001110110 : begin
                   	state <= 10'b0001110111;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001110111 : begin
                   	state <= 10'b0001111000;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001111000 : begin
                   	state <= 10'b0001111001;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hF;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h16;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001111001 : begin
                   	state <= 10'b0001111010;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h16;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001111010 : begin
                   	state <= 10'b0001111011;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h14;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001111011 : begin
                   	state <= 10'b0001111100;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h14;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001111100 : begin
                   	state <= 10'b0001111101;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h11;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h13;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001111101 : begin
                   	state <= 10'b0001111110;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h13;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0001111110 : begin
                   	state <= 10'b0001111111;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0001111111 : begin
                   	state <= 10'b0010000000;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1C;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000000 : begin
                   	state <= 10'b0010000001;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1C;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000001 : begin
                   	state <= 10'b0010000010;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h15;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b0010000010 : begin
                   	state <= 10'b0010000011;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h15;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000011 : begin
                   	state <= 10'b0010000100;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000100 : begin
                   	state <= 10'b0010000101;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1B;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000101 : begin
                   	state <= 10'b0010000110;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1B;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000110 : begin
                   	state <= 10'b0010000111;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010000111 : begin
                   	state <= 10'b0010001000;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001000 : begin
                   	state <= 10'b0010001001;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'hF;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h16;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001001 : begin
                   	state <= 10'b0010001010;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h16;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001010 : begin
                   	state <= 10'b0010001011;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h14;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001011 : begin
                   	state <= 10'b0010001100;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h14;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001100 : begin
                   	state <= 10'b0010001101;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h11;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h13;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001101 : begin
                   	state <= 10'b0010001110;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h13;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001110 : begin
                   	state <= 10'b0010001111;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010001111 : begin
                   	state <= 10'b0010010000;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1C;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010000 : begin
                   	state <= 10'b0010010001;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1C;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010001 : begin
                   	state <= 10'b0010010010;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h15;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010010 : begin
                   	state <= 10'b0010010011;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h15;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010011 : begin
                   	state <= 10'b0010010100;
                   	MultConst_const <= 8'h9;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1B;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010100 : begin
                   	state <= 10'b0010010101;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1B;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010101 : begin
                   	state <= 10'b0010010110;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010110 : begin
                   	state <= 10'b0010010111;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010010111 : begin
                   	state <= 10'b0010011000;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011000 : begin
                   	state <= 10'b0010011001;
                   	MultConst_const <= 8'h2;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'hF;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h16;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011001 : begin
                   	state <= 10'b0010011010;
                   	MultConst_const <= 8'h3;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h16;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'hF;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h14;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011010 : begin
                   	state <= 10'b0010011011;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h14;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011011 : begin
                   	state <= 10'b0010011100;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011100 : begin
                   	state <= 10'b0010011101;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h11;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h13;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011101 : begin
                   	state <= 10'b0010011110;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h13;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011110 : begin
                   	state <= 10'b0010011111;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010011111 : begin
                   	state <= 10'b0010100000;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1C;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100000 : begin
                   	state <= 10'b0010100001;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1C;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100001 : begin
                   	state <= 10'b0010100010;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'hE;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h1B;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100010 : begin
                   	state <= 10'b0010100011;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1B;
                   	MultConst_addr_w <= 5'hB;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h15;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100011 : begin
                   	state <= 10'b0010100100;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h15;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'hB;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100100 : begin
                   	state <= 10'b0010100101;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'hB;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100101 : begin
                   	state <= 10'b0010100110;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'hB;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100110 : begin
                   	state <= 10'b0010100111;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'hB;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010100111 : begin
                   	state <= 10'b0010101000;
                   	MultConst_const <= 8'h25;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hF;
                   	Add_Z__addr_r <= 5'hB;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h16;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101000 : begin
                   	state <= 10'b0010101001;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h16;
                   	MultConst_addr_w <= 5'hB;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101001 : begin
                   	state <= 10'b0010101010;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'hB;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h14;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101010 : begin
                   	state <= 10'b0010101011;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h14;
                   	MultConst_addr_w <= 5'hB;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101011 : begin
                   	state <= 10'b0010101100;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h11;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'hB;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h13;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h14;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101100 : begin
                   	state <= 10'b0010101101;
                   	MultConst_const <= 8'h2;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h13;
                   	MultConst_addr_w <= 5'hB;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'hD;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h14;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101101 : begin
                   	state <= 10'b0010101110;
                   	MultConst_const <= 8'h3;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101110 : begin
                   	state <= 10'b0010101111;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1C;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010101111 : begin
                   	state <= 10'b0010110000;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1C;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110000 : begin
                   	state <= 10'b0010110001;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h15;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110001 : begin
                   	state <= 10'b0010110010;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h15;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110010 : begin
                   	state <= 10'b0010110011;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1B;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110011 : begin
                   	state <= 10'b0010110100;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1B;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'hC;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1B;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110100 : begin
                   	state <= 10'b0010110101;
                   	MultConst_const <= 8'h2;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'hE;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'hB;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1B;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110101 : begin
                   	state <= 10'b0010110110;
                   	MultConst_const <= 8'h3;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h2;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110110 : begin
                   	state <= 10'b0010110111;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h16;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010110111 : begin
                   	state <= 10'b0010111000;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h16;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h13;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111000 : begin
                   	state <= 10'b0010111001;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h13;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111001 : begin
                   	state <= 10'b0010111010;
                   	MultConst_const <= 8'hf4;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111010 : begin
                   	state <= 10'b0010111011;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h11;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111011 : begin
                   	state <= 10'b0010111100;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111100 : begin
                   	state <= 10'b0010111101;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h9;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111101 : begin
                   	state <= 10'b0010111110;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1C;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111110 : begin
                   	state <= 10'b0010111111;
                   	MultConst_const <= 8'h2;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1C;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h8;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0010111111 : begin
                   	state <= 10'b0011000000;
                   	MultConst_const <= 8'h3;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'hF;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h15;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000000 : begin
                   	state <= 10'b0011000001;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h15;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000001 : begin
                   	state <= 10'b0011000010;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000010 : begin
                   	state <= 10'b0011000011;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h16;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000011 : begin
                   	state <= 10'b0011000100;
                   	MultConst_const <= 8'h2;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h16;
                   	MultConst_addr_w <= 5'h8;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000100 : begin
                   	state <= 10'b0011000101;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000101 : begin
                   	state <= 10'b0011000110;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h9;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h5;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000110 : begin
                   	state <= 10'b0011000111;
                   	MultConst_const <= 8'h2;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h11;
                   	MultConst_addr_w <= 5'h11;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'hE;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011000111 : begin
                   	state <= 10'b0011001000;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h4;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001000 : begin
                   	state <= 10'b0011001001;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h9;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h13;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001001 : begin
                   	state <= 10'b0011001010;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h13;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001010 : begin
                   	state <= 10'b0011001011;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h9;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h1C;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h13;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001011 : begin
                   	state <= 10'b0011001100;
                   	MultConst_const <= 8'h2;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1C;
                   	MultConst_addr_w <= 5'hD;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h13;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001100 : begin
                   	state <= 10'b0011001101;
                   	MultConst_const <= 8'h3;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hC;
                   	MultConst_addr_w <= 5'h11;
                   	Square_addr_w <= 5'h6;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Add_Z__addr_r <= 5'hE;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001101 : begin
                   	state <= 10'b0011001110;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001110 : begin
                   	state <= 10'b0011001111;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'h10;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h2;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h15;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011001111 : begin
                   	state <= 10'b0011010000;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h15;
                   	MultConst_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h9;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011010000 : begin
                   	state <= 10'b0011010001;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'h9;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011010001 : begin
                   	state <= 10'b0011010010;
                   	MultConst_const <= 8'h2;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'h5;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h16;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011010010 : begin
                   	state <= 10'b0011010011;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h16;
                   	MultConst_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011010011 : begin
                   	state <= 10'b0011010100;
                   	MultConst_const <= 8'hb5;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'hE;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011010100 : begin
                   	state <= 10'b0011010101;
                   	MultConst_const <= 8'hb5;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h9;
                   	MultConst_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'h1B;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011010101 : begin
                   	state <= 10'b0011010110;
                   	MultConst_const <= 8'h2;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'h12;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011010110 : begin
                   	state <= 10'b0011010111;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h11;
                   	MultConst_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'h9;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b0011010111 : begin
                   	state <= 10'b0011011000;
                   	MultConst_const <= 8'hb5;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h2;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h16;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011000 : begin
                   	state <= 10'b0011011001;
                   	MultConst_const <= 8'h2;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1D;
                   	MultConst_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h8;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h16;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h16;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011001 : begin
                   	state <= 10'b0011011010;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h8;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h16;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011010 : begin
                   	state <= 10'b0011011011;
                   	MultConst_const <= 8'h2;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h16;
                   	MultConst_addr_w <= 5'h8;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Add_Z__addr_r <= 5'h1B;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011011 : begin
                   	state <= 10'b0011011100;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1B;
                   	MultConst_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1C;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h11;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011100 : begin
                   	state <= 10'b0011011101;
                   	MultConst_const <= 8'h2;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1C;
                   	MultConst_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'hE;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h15;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h11;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011101 : begin
                   	state <= 10'b0011011110;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h15;
                   	MultConst_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'hD;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011110 : begin
                   	state <= 10'b0011011111;
                   	MultConst_const <= 8'h2;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h5;
                   	MultConst_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h13;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011011111 : begin
                   	state <= 10'b0011100000;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h11;
                   	MultConst_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'h9;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1C;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100000 : begin
                   	state <= 10'b0011100001;
                   	MultConst_const <= 8'h2;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h14;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1C;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100001 : begin
                   	state <= 10'b0011100010;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1A;
                   	MultConst_addr_w <= 5'h7;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h15;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100010 : begin
                   	state <= 10'b0011100011;
                   	MultConst_const <= 8'h2;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h15;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100011 : begin
                   	state <= 10'b0011100100;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h18;
                   	MultConst_addr_w <= 5'h5;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Add_Z__addr_r <= 5'h8;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100100 : begin
                   	state <= 10'b0011100101;
                   	MultConst_const <= 8'h2;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h1C;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100101 : begin
                   	state <= 10'b0011100110;
                   	MultConst_const <= 8'h3;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1E;
                   	MultConst_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h12;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1C;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011100110 : begin
                   	state <= 10'b0011100111;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1C;
                   	Add_Z__addr_r <= 5'h11;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h10;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   end
                   10'b0011100111 : begin
                   	state <= 10'b0011101000;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h19;
                   	Add_Z__addr_r <= 5'h15;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101000 : begin
                   	state <= 10'b0011101001;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h17;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Add_Z__addr_r <= 5'h15;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101001 : begin
                   	state <= 10'b0011101010;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h15;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Add_Z__addr_r <= 5'h13;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101010 : begin
                   	state <= 10'b0011101011;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h13;
                   	Add_Z__addr_r <= 5'hD;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h14;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101011 : begin
                   	state <= 10'b0011101100;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h14;
                   	Add_Z__addr_r <= 5'hC;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   end
                   10'b0011101100 : begin
                   	state <= 10'b0011101101;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h12;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h9;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   end
                   10'b0011101101 : begin
                   	state <= 10'b0011101110;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'h8;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101110 : begin
                   	state <= 10'b0011101111;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011101111 : begin
                   	state <= 10'b0011110000;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110000 : begin
                   	state <= 10'b0011110001;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110001 : begin
                   	state <= 10'b0011110010;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110010 : begin
                   	state <= 10'b0011110011;
                   	Add_Z__addr_r <= 5'h5;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h4;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   end
                   10'b0011110011 : begin
                   	state <= 10'b0011110100;
                   	round_pt[6*8*v-1 -: 8*v] <= Add_P;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   end
                   10'b0011110100 : begin
                   	state <= 10'b0011110101;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h1E;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h1D;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110101 : begin
                   	state <= 10'b0011110110;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110110 : begin
                   	state <= 10'b0011110111;
                   	round_pt[9*8*v-1 -: 8*v] <= Add_P;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h1C;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h1B;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011110111 : begin
                   	state <= 10'b0011111000;
                   	Add_Z__addr_r <= 5'h1A;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h19;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111000 : begin
                   	state <= 10'b0011111001;
                   	round_pt[12*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h18;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h17;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111001 : begin
                   	state <= 10'b0011111010;
                   	round_pt[5*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h16;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h15;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111010 : begin
                   	state <= 10'b0011111011;
                   	round_pt[15*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h14;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h13;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111011 : begin
                   	state <= 10'b0011111100;
                   	round_pt[16*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h12;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h11;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111100 : begin
                   	state <= 10'b0011111101;
                   	round_pt[8*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111101 : begin
                   	state <= 10'b0011111110;
                   	round_pt[7*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'hE;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'hD;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111110 : begin
                   	state <= 10'b0011111111;
                   	round_pt[11*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'hC;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0011111111 : begin
                   	state <= 10'b0100000000;
                   	round_pt[2*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h9;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0100000000 : begin
                   	state <= 10'b0100000001;
                   	round_pt[3*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h8;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0100000001 : begin
                   	state <= 10'b0100000010;
                   	round_pt[10*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0100000010 : begin
                   	state <= 10'b0100000011;
                   	round_pt[14*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0100000011 : begin
                   	state <= 10'b0100000100;
                   	round_pt[13*8*v-1 -: 8*v] <= Add_P;
                   	round_count <= round_count + 1; // sen_ding this two cycles early to receive values from ks earlier
                   	Add_Z__addr_r <= 5'h2;
                   	Add_Z__addr_r_BRAM <= BRAM_add;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b0100000100 : begin
                   	state <= 10'b0100000101;
                   	round_pt[1*8*v-1 -: 8*v] <= Add_P;
                   end
                   10'b0100000101 : begin
                   	state <= {is_last, 9'b000000000};
                   	round_pt[4*8*v-1 -: 8*v] <= Add_P;
                   end
                   // LAST ROUND STARTS HERE
                   10'b1000000000 : begin
                   	state <= 10'b1000000001;
                   	Add_Z_addr_r <= 5'h10; // addr of byte F
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h10; // addr of byte F
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   end
                   10'b1000000001 : begin
                   	state <= 10'b1000000010;
                   	Add_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hF; // addr of byte E
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hF; // addr of byte E
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h5;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000000010 : begin
                   	state <= 10'b1000000011;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hE; // addr of byte D
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hE; // addr of byte D
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h8;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h5;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000000011 : begin
                   	state <= 10'b1000000100;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hD; // addr of byte C
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hD; // addr of byte C
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h10;
                   	Mult_addr_w <= 5'h15;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h8;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h15;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000000100 : begin
                   	state <= 10'b1000000101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hC; // addr of byte B
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hC; // addr of byte B
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h4;
                   	Mult_addr_w <= 5'h19;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h5;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000000101 : begin
                   	state <= 10'b1000000110;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hB; // addr of byte A
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hB; // addr of byte A
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h5;
                   	Mult_addr_w <= 5'h16;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h10;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000000110 : begin
                   	state <= 10'b1000000111;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'hA; // addr of byte 9
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'hA; // addr of byte 9
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h6;
                   	Mult_addr_w <= 5'h8;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h15;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h19;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000000111 : begin
                   	state <= 10'b1000001000;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h9; // addr of byte 8
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h9; // addr of byte 8
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h7;
                   	Mult_addr_w <= 5'h15;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h8;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000001000 : begin
                   	state <= 10'b1000001001;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h8; // addr of byte 7
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h8; // addr of byte 7
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h8;
                   	Mult_addr_w <= 5'h13;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h4;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000001001 : begin
                   	state <= 10'b1000001010;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h7; // addr of byte 6
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h7; // addr of byte 6
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h9;
                   	Mult_addr_w <= 5'h9;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h5;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000001010 : begin
                   	state <= 10'b1000001011;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h6; // addr of byte 5
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h6; // addr of byte 5
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hA;
                   	Mult_addr_w <= 5'h1C;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h10;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000001011 : begin
                   	state <= 10'b1000001100;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h5; // addr of byte 4
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h5; // addr of byte 4
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h10;
                   	Mult_addr_w <= 5'hE;
                   	Square_addr_w <= 5'h3;
                   	Mult_Z_addr_r <= 5'h3;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h6;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h15;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000001100 : begin
                   	state <= 10'b1000001101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h4; // addr of byte 3
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h4; // addr of byte 3
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hB;
                   	Mult_addr_w <= 5'h15;
                   	Square_addr_w <= 5'h3;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000001101 : begin
                   	state <= 10'b1000001110;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h3; // addr of byte 2
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h3; // addr of byte 2
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hC;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h19;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000001110 : begin
                   	state <= 10'b1000001111;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h2; // addr of byte 1
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h2; // addr of byte 1
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hD;
                   	Mult_addr_w <= 5'h19;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h7;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000001111 : begin
                   	state <= 10'b1000010000;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z_addr_r <= 5'h1; // addr of byte 0
                   	Add_Z_addr_r_BRAM <= BRAM_PT; // take from plaintext
                   	Add_Z__addr_r <= 5'h1; // addr of byte 0
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hE;
                   	Mult_addr_w <= 5'h12;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h8;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000010000 : begin
                   	state <= 10'b1000010001;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	Mult_addr_w <= 5'h18;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h4;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000010001 : begin
                   	state <= 10'b1000010010;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h10;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h9;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000010010 : begin
                   	state <= 10'b1000010011;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h17;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h8;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h1C;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000010011 : begin
                   	state <= 10'b1000010100;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h8;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h5;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000010100 : begin
                   	state <= 10'b1000010101;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hC;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hA;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000010101 : begin
                   	state <= 10'b1000010110;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h1B;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h10;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000010110 : begin
                   	state <= 10'b1000010111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h1A;
                   	Square_addr_w <= 5'h3;
                   	Square_Z_addr_r <= 5'h15;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000010111 : begin
                   	state <= 10'b1000011000;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h6;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000011000 : begin
                   	state <= 10'b1000011001;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h7;
                   	Square_addr_w <= 5'hA;
                   	Mult_Z_addr_r <= 5'hA;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hB;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000011001 : begin
                   	state <= 10'b1000011010;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h14;
                   	Square_addr_w <= 5'hA;
                   	Mult_Z_addr_r <= 5'hA;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hC;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h19;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000011010 : begin
                   	state <= 10'b1000011011;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h19;
                   	Square_addr_w <= 5'hA;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000011011 : begin
                   	state <= 10'b1000011100;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hD;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h12;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000011100 : begin
                   	state <= 10'b1000011101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h11;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h7;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000011101 : begin
                   	state <= 10'b1000011110;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hE;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000011110 : begin
                   	state <= 10'b1000011111;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hD;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h9;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h18;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000011111 : begin
                   	state <= 10'b1000100000;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h9;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h8;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1000100000 : begin
                   	state <= 10'b1000100001;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h2;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hF;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h17;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000100001 : begin
                   	state <= 10'b1000100010;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hF;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h9;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000100010 : begin
                   	state <= 10'b1000100011;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h8;
                   	Square_addr_w <= 5'hB;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000100011 : begin
                   	state <= 10'b1000100100;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1C;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h1B;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000100100 : begin
                   	state <= 10'b1000100101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h1C;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hA;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000100101 : begin
                   	state <= 10'b1000100110;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hB;
                   	Square_addr_w <= 5'h3;
                   	Mult_Z_addr_r <= 5'h3;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h16;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h1A;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000100110 : begin
                   	state <= 10'b1000100111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h16;
                   	Square_addr_w <= 5'h3;
                   	Mult_Z_addr_r <= 5'h3;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h10;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h16;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000100111 : begin
                   	state <= 10'b1000101000;
                   	MultConst_const <= 8'h8f;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	can_supply_last <= 1'b1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Mult_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hF;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h15;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h14;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000101000 : begin
                   	state <= 10'b1000101001;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h10;
                   	Mult_addr_w <= 5'h15;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hB;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000101001 : begin
                   	state <= 10'b1000101010;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h5;
                   	Square_addr_w <= 5'hA;
                   	Square_Z_addr_r <= 5'h19;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000101010 : begin
                   	state <= 10'b1000101011;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hD;
                   	Mult_Z_addr_r <= 5'hD;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hC;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000101011 : begin
                   	state <= 10'b1000101100;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h4;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h12;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h11;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000101100 : begin
                   	state <= 10'b1000101101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h12;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hD;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000101101 : begin
                   	state <= 10'b1000101110;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h4;
                   	Mult_Z_addr_r <= 5'h4;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hE;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000101110 : begin
                   	state <= 10'b1000101111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h9;
                   	Square_addr_w <= 5'h9;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000101111 : begin
                   	state <= 10'b1000110000;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h2;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h18;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000110000 : begin
                   	state <= 10'b1000110001;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h18;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h17;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000110001 : begin
                   	state <= 10'b1000110010;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h17;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hF;
                   	Mult_Z__addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000110010 : begin
                   	state <= 10'b1000110011;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h1;
                   	Square_addr_w <= 5'hB;
                   	Square_Z_addr_r <= 5'h1C;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000110011 : begin
                   	state <= 10'b1000110100;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h2;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000110100 : begin
                   	state <= 10'b1000110101;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h10;
                   	Mult_Z_addr_r <= 5'h10;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1B;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h16;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000110101 : begin
                   	state <= 10'b1000110110;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h16;
                   	Square_addr_w <= 5'h10;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000110110 : begin
                   	state <= 10'b1000110111;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h10;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'h3;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1A;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h15;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000110111 : begin
                   	state <= 10'b1000111000;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h10;
                   	Mult_addr_w <= 5'h15;
                   	Square_addr_w <= 5'h3;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111000 : begin
                   	state <= 10'b1000111001;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hF;
                   	Mult_Z_addr_r <= 5'hF;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h14;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111001 : begin
                   	state <= 10'b1000111010;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h14;
                   	Square_addr_w <= 5'hA;
                   	Mult_Z_addr_r <= 5'hA;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h13;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111010 : begin
                   	state <= 10'b1000111011;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h13;
                   	Square_addr_w <= 5'hD;
                   	Mult_Z_addr_r <= 5'hD;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h19;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h13;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h12;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000111011 : begin
                   	state <= 10'b1000111100;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Mult_addr_w <= 5'h12;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hD;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111100 : begin
                   	state <= 10'b1000111101;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h11;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111101 : begin
                   	state <= 10'b1000111110;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h11;
                   	Square_addr_w <= 5'h4;
                   	Mult_Z_addr_r <= 5'h4;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hD;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1000111110 : begin
                   	state <= 10'b1000111111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hD;
                   	Square_addr_w <= 5'h9;
                   	Square_Z_addr_r <= 5'h18;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1000111111 : begin
                   	state <= 10'b1001000000;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h4;
                   	Square_Z_addr_r <= 5'h17;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001000000 : begin
                   	state <= 10'b1001000001;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hC;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001000001 : begin
                   	state <= 10'b1001000010;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h5;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hF;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001000010 : begin
                   	state <= 10'b1001000011;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hF;
                   	Square_addr_w <= 5'hB;
                   	Mult_Z_addr_r <= 5'hB;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hE;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001000011 : begin
                   	state <= 10'b1001000100;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hE;
                   	Square_addr_w <= 5'h2;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001000100 : begin
                   	state <= 10'b1001000101;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h10;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h16;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001000101 : begin
                   	state <= 10'b1001000110;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h10;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001000110 : begin
                   	state <= 10'b1001000111;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h10;
                   	Square_addr_w <= 5'h3;
                   	Square_Z_addr_r <= 5'h15;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001000111 : begin
                   	state <= 10'b1001001000;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h5;
                   	Square_Z_addr_r <= 5'h14;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001001000 : begin
                   	state <= 10'b1001001001;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hA;
                   	Square_Z_addr_r <= 5'h13;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001001001 : begin
                   	state <= 10'b1001001010;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hF;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001001010 : begin
                   	state <= 10'b1001001011;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h12;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001001011 : begin
                   	state <= 10'b1001001100;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	Square_addr_w <= 5'h6;
                   	Square_Z_addr_r <= 5'h11;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001001100 : begin
                   	state <= 10'b1001001101;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h8;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001001101 : begin
                   	state <= 10'b1001001110;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h9;
                   	Mult_Z_addr_r <= 5'h9;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h10;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001001110 : begin
                   	state <= 10'b1001001111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Mult_addr_w <= 5'hD;
                   	Square_addr_w <= 5'h9;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001001111 : begin
                   	state <= 10'b1001010000;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h4;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010000 : begin
                   	state <= 10'b1001010001;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hD;
                   	Square_addr_w <= 5'hC;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001010001 : begin
                   	state <= 10'b1001010010;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'h7;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001010010 : begin
                   	state <= 10'b1001010011;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hE;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010011 : begin
                   	state <= 10'b1001010100;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'h2;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hC;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010100 : begin
                   	state <= 10'b1001010101;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	Mult_addr_w <= 5'hC;
                   	Square_addr_w <= 5'h10;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010101 : begin
                   	state <= 10'b1001010110;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h10;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010110 : begin
                   	state <= 10'b1001010111;
                   	MultConst_const <= 8'h8f;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'h10;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h3;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Mult_Z_addr_r <= 5'h3;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h7;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001010111 : begin
                   	state <= 10'b1001011000;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hC;
                   	Mult_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h5;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011000 : begin
                   	state <= 10'b1001011001;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hA;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011001 : begin
                   	state <= 10'b1001011010;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	Square_addr_w <= 5'hF;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011010 : begin
                   	state <= 10'b1001011011;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'hD;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hA;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011011 : begin
                   	state <= 10'b1001011100;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	Mult_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h6;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011100 : begin
                   	state <= 10'b1001011101;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h8;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001011101 : begin
                   	state <= 10'b1001011110;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	Square_addr_w <= 5'hD;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011110 : begin
                   	state <= 10'b1001011111;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hD;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001011111 : begin
                   	state <= 10'b1001100000;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'hD;
                   	Square_addr_w <= 5'h4;
                   	Mult_Z_addr_r <= 5'h4;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h2;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100000 : begin
                   	state <= 10'b1001100001;
                   	Mult_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Mult_addr_w <= 5'h2;
                   	Square_addr_w <= 5'hC;
                   	Mult_Z_addr_r <= 5'hC;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h8;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100001 : begin
                   	state <= 10'b1001100010;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Mult_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h7;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100010 : begin
                   	state <= 10'b1001100011;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'h9;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hE;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100011 : begin
                   	state <= 10'b1001100100;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001100100 : begin
                   	state <= 10'b1001100101;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h10;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100101 : begin
                   	state <= 10'b1001100110;
                   	MultConst_const <= 8'h5;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h10;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hC;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'hB;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'hB;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001100110 : begin
                   	state <= 10'b1001100111;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hC;
                   	Mult_addr_w <= 5'h7;
                   	Square_addr_w <= 5'hB;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001100111 : begin
                   	state <= 10'b1001101000;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'h5;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h6;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101000 : begin
                   	state <= 10'b1001101001;
                   	MultConst_const <= 8'h8f;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'hB;
                   	Mult_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hA;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Mult_Z_addr_r <= 5'hA;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h5;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101001 : begin
                   	state <= 10'b1001101010;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'h7;
                   	Mult_addr_w <= 5'h5;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hF;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001101010 : begin
                   	state <= 10'b1001101011;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101011 : begin
                   	state <= 10'b1001101100;
                   	MultConst_const <= 8'h8f;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h6;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Mult_Z_addr_r <= 5'h6;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h4;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101100 : begin
                   	state <= 10'b1001101101;
                   	MultConst_const <= 8'h5;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h5;
                   	Mult_addr_w <= 5'h4;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'h8;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h3;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101101 : begin
                   	state <= 10'b1001101110;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'hA;
                   	Mult_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hD;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001101110 : begin
                   	state <= 10'b1001101111;
                   	MultConst_const <= 8'h9;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h4;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hD;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Mult_Z_addr_r <= 5'h9;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h9;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001101111 : begin
                   	state <= 10'b1001110000;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'hD;
                   	Mult_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h9;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001110000 : begin
                   	state <= 10'b1001110001;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h9;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001110001 : begin
                   	state <= 10'b1001110010;
                   	MultConst_const <= 8'h8f;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'h9;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h7;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	Mult_Z_addr_r <= 5'h7;
                   	Mult_Z_addr_r_BRAM <= BRAM_sq;
                   	Mult_Z__addr_r <= 5'h1;
                   	Mult_Z__addr_r_BRAM <= BRAM_mul;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001110010 : begin
                   	state <= 10'b1001110011;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Mult_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	Mult_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001110011 : begin
                   	state <= 10'b1001110100;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_mul;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001110100 : begin
                   	state <= 10'b1001110101;
                   	MultConst_const <= 8'h8f;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r_BRAM <= BRAM_mask; // take from Mask
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hC;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_mc;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001110101 : begin
                   	state <= 10'b1001110110;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h10;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001110110 : begin
                   	state <= 10'b1001110111;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h10;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hC;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001110111 : begin
                   	state <= 10'b1001111000;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hC;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001111000 : begin
                   	state <= 10'b1001111001;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hF;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001111001 : begin
                   	state <= 10'b1001111010;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001111010 : begin
                   	state <= 10'b1001111011;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001111011 : begin
                   	state <= 10'b1001111100;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001111100 : begin
                   	state <= 10'b1001111101;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h5;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001111101 : begin
                   	state <= 10'b1001111110;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h4;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1001111110 : begin
                   	state <= 10'b1001111111;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h4;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hD;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1001111111 : begin
                   	state <= 10'b1010000000;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hD;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000000 : begin
                   	state <= 10'b1010000001;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h9;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000001 : begin
                   	state <= 10'b1010000010;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h9;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_mul;
                   end
                   10'b1010000010 : begin
                   	state <= 10'b1010000011;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000011 : begin
                   	state <= 10'b1010000100;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'h10;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h10;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000100 : begin
                   	state <= 10'b1010000101;
                   	MultConst_const <= 8'h5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h10;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000101 : begin
                   	state <= 10'b1010000110;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000110 : begin
                   	state <= 10'b1010000111;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hC;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010000111 : begin
                   	state <= 10'b1010001000;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hC;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001000 : begin
                   	state <= 10'b1010001001;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'hF;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001001 : begin
                   	state <= 10'b1010001010;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001010 : begin
                   	state <= 10'b1010001011;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001011 : begin
                   	state <= 10'b1010001100;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001100 : begin
                   	state <= 10'b1010001101;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h5;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001101 : begin
                   	state <= 10'b1010001110;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h4;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001110 : begin
                   	state <= 10'b1010001111;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h4;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hD;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010001111 : begin
                   	state <= 10'b1010010000;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hD;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010000 : begin
                   	state <= 10'b1010010001;
                   	MultConst_const <= 8'h9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h9;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010001 : begin
                   	state <= 10'b1010010010;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h9;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010010 : begin
                   	state <= 10'b1010010011;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h10;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010011 : begin
                   	state <= 10'b1010010100;
                   	MultConst_const <= 8'h9;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h10;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h10;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010100 : begin
                   	state <= 10'b1010010101;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010101 : begin
                   	state <= 10'b1010010110;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h10;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010110 : begin
                   	state <= 10'b1010010111;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h10;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hC;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010010111 : begin
                   	state <= 10'b1010011000;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r <= 5'h4; // addr of byte 3
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hC;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h6;
                   	Add_Z_addr_r <= 5'h10;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011000 : begin
                   	state <= 10'b1010011001;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'hF;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011001 : begin
                   	state <= 10'b1010011010;
                   	round_pt[4*8*v-1 -: 8*v] <= Add_P;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011010 : begin
                   	state <= 10'b1010011011;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'hF;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011011 : begin
                   	state <= 10'b1010011100;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011100 : begin
                   	state <= 10'b1010011101;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011101 : begin
                   	state <= 10'b1010011110;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h5;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011110 : begin
                   	state <= 10'b1010011111;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h4;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010011111 : begin
                   	state <= 10'b1010100000;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h4;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hD;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100000 : begin
                   	state <= 10'b1010100001;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hD;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100001 : begin
                   	state <= 10'b1010100010;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h9;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100010 : begin
                   	state <= 10'b1010100011;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h9;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100011 : begin
                   	state <= 10'b1010100100;
                   	MultConst_const <= 8'hf9;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'hE;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100100 : begin
                   	state <= 10'b1010100101;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100101 : begin
                   	state <= 10'b1010100110;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100110 : begin
                   	state <= 10'b1010100111;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hC;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hF;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010100111 : begin
                   	state <= 10'b1010101000;
                   	MultConst_const <= 8'h25;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'hC;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'hF;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hF;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101000 : begin
                   	state <= 10'b1010101001;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101001 : begin
                   	state <= 10'b1010101010;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101010 : begin
                   	state <= 10'b1010101011;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101011 : begin
                   	state <= 10'b1010101100;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hF;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101100 : begin
                   	state <= 10'b1010101101;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h5;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101101 : begin
                   	state <= 10'b1010101110;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_Z__addr_r <= 5'h7; // addr of byte 6
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hA;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h9;
                   	Add_Z_addr_r <= 5'hF;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101110 : begin
                   	state <= 10'b1010101111;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'hD;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'hD;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010101111 : begin
                   	state <= 10'b1010110000;
                   	round_pt[7*8*v-1 -: 8*v] <= Add_P;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hD;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h4;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hE;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110000 : begin
                   	state <= 10'b1010110001;
                   	MultConst_const <= 8'hf4;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h4;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'hE;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hE;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110001 : begin
                   	state <= 10'b1010110010;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h9;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110010 : begin
                   	state <= 10'b1010110011;
                   	MultConst_const <= 8'h25;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h9;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110011 : begin
                   	state <= 10'b1010110100;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110100 : begin
                   	state <= 10'b1010110101;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110101 : begin
                   	state <= 10'b1010110110;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hE;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'hC;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'hC;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110110 : begin
                   	state <= 10'b1010110111;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'hC;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010110111 : begin
                   	state <= 10'b1010111000;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'hB;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111000 : begin
                   	state <= 10'b1010111001;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_Z__addr_r <= 5'hA; // addr of byte 9
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'hB;
                   	Square_addr_w <= 5'h4;
                   	Add_Z_addr_r <= 5'hE;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hD;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111001 : begin
                   	state <= 10'b1010111010;
                   	MultConst_const <= 8'hf4;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'hD;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hD;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111010 : begin
                   	state <= 10'b1010111011;
                   	round_pt[10*8*v-1 -: 8*v] <= Add_P;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111011 : begin
                   	state <= 10'b1010111100;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h6;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'hA;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111100 : begin
                   	state <= 10'b1010111101;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111101 : begin
                   	state <= 10'b1010111110;
                   	MultConst_const <= 8'hf4;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h5;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h4;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111110 : begin
                   	state <= 10'b1010111111;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hD;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h1;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hC;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1010111111 : begin
                   	state <= 10'b1011000000;
                   	MultConst_const <= 8'hf4;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'hD;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'hC;
                   	Add_Z__addr_r <= 5'h9;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h9;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hC;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'hB;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000000 : begin
                   	state <= 10'b1011000001;
                   	MultConst_const <= 8'hb5;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h9;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'hB;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hB;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000001 : begin
                   	state <= 10'b1011000010;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'h8;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000010 : begin
                   	state <= 10'b1011000011;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	Square_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000011 : begin
                   	state <= 10'b1011000100;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_Z__addr_r <= 5'hD; // addr of byte C
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h2;
                   	Square_addr_w <= 5'h5;
                   	Add_Z_addr_r <= 5'hD;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'hA;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000100 : begin
                   	state <= 10'b1011000101;
                   	Square_BRAM_en <= 1;
                   	Square_addr_w <= 5'hA;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'hA;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000101 : begin
                   	state <= 10'b1011000110;
                   	round_pt[13*8*v-1 -: 8*v] <= Add_P;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h1;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h4;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hC;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000110 : begin
                   	state <= 10'b1011000111;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'hC;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h9;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011000111 : begin
                   	state <= 10'b1011001000;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'hB;
                   	Square_addr_w <= 5'h9;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h9;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001000 : begin
                   	state <= 10'b1011001001;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h8;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001001 : begin
                   	state <= 10'b1011001010;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h8;
                   	Add_Z__addr_r <= 5'h5;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h8;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001010 : begin
                   	state <= 10'b1011001011;
                   	MultConst_const <= 8'hb5;
                   	Square_BRAM_en <= 1;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h5;
                   	MultConst_addr_w <= 5'h1;
                   	Square_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	Square_Z_addr_r <= 5'h7;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001011 : begin
                   	state <= 10'b1011001100;
                   	Add_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'hA;
                   	Square_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h4;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h7;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h6;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001100 : begin
                   	state <= 10'b1011001101;
                   	MultConst_const <= 8'hb5;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z__addr_r <= 5'h10; // addr of byte F
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h4;
                   	MultConst_addr_w <= 5'h7;
                   	Square_addr_w <= 5'h6;
                   	Add_Z_addr_r <= 5'hC;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h6;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h5;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001101 : begin
                   	state <= 10'b1011001110;
                   	MultConst_const <= 8'hb5;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h6;
                   	Square_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h5;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h4;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001110 : begin
                   	state <= 10'b1011001111;
                   	round_pt[16*8*v-1 -: 8*v] <= Add_P;
                   	MultConst_const <= 8'hb5;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_Z__addr_r <= 5'h3; // addr of byte 2
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h3;
                   	MultConst_addr_w <= 5'h5;
                   	Square_addr_w <= 5'h4;
                   	Add_Z_addr_r <= 5'hB;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h4;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h3;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011001111 : begin
                   	state <= 10'b1011010000;
                   	MultConst_const <= 8'hb5;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	MultConst_addr_w <= 5'h4;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h9;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h2;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011010000 : begin
                   	state <= 10'b1011010001;
                   	round_pt[3*8*v-1 -: 8*v] <= Add_P;
                   	MultConst_const <= 8'hb5;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h9;
                   	MultConst_addr_w <= 5'h3;
                   	Square_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h2;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h3;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   	Square_Z_addr_r <= 5'h1;
                   	Square_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011010001 : begin
                   	state <= 10'b1011010010;
                   	MultConst_const <= 8'hb5;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Square_BRAM_en <= 1;
                   	Add_addr_w <= 5'h2;
                   	MultConst_addr_w <= 5'h2;
                   	Square_addr_w <= 5'h2;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   	MultConst_Z_addr_r <= 5'h2;
                   	MultConst_Z_addr_r_BRAM <= BRAM_sq;
                   end
                   10'b1011010010 : begin
                   	state <= 10'b1011010011;
                   	MultConst_const <= 8'hb5;
                   	Add_BRAM_en <= 1;
                   	MultConst_BRAM_en <= 1;
                   	Add_addr_w <= 5'h8;
                   	MultConst_addr_w <= 5'h1;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_sq;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011010011 : begin
                   	state <= 10'b1011010100;
                   	Add_BRAM_en <= 1;
                   	Add_Z__addr_r <= 5'h6; // addr of byte 5
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h1;
                   	Add_Z_addr_r <= 5'hA;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011010100 : begin
                   	state <= 10'b1011010101;
                   	Add_Z__addr_r <= 5'h7;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011010101 : begin
                   	state <= 10'b1011010110;
                   	round_pt[6*8*v-1 -: 8*v] <= Add_P;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h7;
                   	Add_Z__addr_r <= 5'h6;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011010110 : begin
                   	state <= 10'b1011010111;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h6;
                   	Add_Z__addr_r <= 5'h5;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011010111 : begin
                   	state <= 10'b1011011000;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h5;
                   	Add_Z__addr_r <= 5'h4;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h4;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011000 : begin
                   	state <= 10'b1011011001;
                   	Add_BRAM_en <= 1;
                   	Add_Z__addr_r <= 5'h9; // addr of byte 8
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h4;
                   	Add_Z_addr_r <= 5'h9;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011001 : begin
                   	state <= 10'b1011011010;
                   	Add_Z__addr_r <= 5'h3;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011010 : begin
                   	state <= 10'b1011011011;
                   	round_pt[9*8*v-1 -: 8*v] <= Add_P;
                   	Add_BRAM_en <= 1;
                   	Add_addr_w <= 5'h3;
                   	Add_Z__addr_r <= 5'h2;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011011 : begin
                   	state <= 10'b1011011100;
                   	Add_BRAM_en <= 1;
                   	Add_Z__addr_r <= 5'hC; // addr of byte B
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h2;
                   	Add_Z_addr_r <= 5'h8;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011100 : begin
                   	state <= 10'b1011011101;
                   	Add_Z__addr_r <= 5'h1;
                   	Add_Z__addr_r_BRAM <= BRAM_mc;
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011101 : begin
                   	state <= 10'b1011011110;
                   	round_pt[12*8*v-1 -: 8*v] <= Add_P;
                   	Add_BRAM_en <= 1;
                   	Add_Z__addr_r <= 5'hF; // addr of byte E
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_addr_w <= 5'h1;
                   	Add_Z_addr_r <= 5'h7;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011110 : begin
                   	state <= 10'b1011011111;
                   	Add_Z__addr_r <= 5'h2; // addr of byte 1
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_Z_addr_r <= 5'h6;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011011111 : begin
                   	state <= 10'b1011100000;
                   	round_pt[15*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h5; // addr of byte 4
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_Z_addr_r <= 5'h5;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011100000 : begin
                   	state <= 10'b1011100001;
                   	round_pt[2*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h8; // addr of byte 7
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_Z_addr_r <= 5'h4;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011100001 : begin
                   	state <= 10'b1011100010;
                   	round_pt[5*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'hB; // addr of byte A
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_Z_addr_r <= 5'h3;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011100010 : begin
                   	state <= 10'b1011100011;
                   	round_pt[8*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'hE; // addr of byte D
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_Z_addr_r <= 5'h2;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011100011 : begin
                   	state <= 10'b1011100100;
                   	round_pt[11*8*v-1 -: 8*v] <= Add_P;
                   	Add_Z__addr_r <= 5'h1; // addr of byte 0
                   	Add_Z__addr_r_BRAM <= BRAM_KS; // take from key
                   	Add_Z_addr_r <= 5'h1;
                   	Add_Z_addr_r_BRAM <= BRAM_add;
                   end
                   10'b1011100100 : begin
                   	state <= 10'b1011100101;
                   	round_pt[14*8*v-1 -: 8*v] <= Add_P;
                   end
                   10'b1011100101 : begin
                   	state <= 10'b1111111100;
                   	round_pt[1*8*v-1 -: 8*v] <= Add_P;
                   	is_busy <= 1'b0;
                   end
                   default : begin
                   	state <= 10'b1111111100;
                   end
                endcase
            end
        end
    end


endmodule